//: version "1.8.7"

module OR(n, p, R, B, A, z);
//: interface  /sz:(40, 40) /bd:[ ]
output p;    //: /sn:0 /dp:1 {0}(627,247)(659,247){1}
output z;    //: /sn:0 /dp:1 {0}(572,286)(593,286){1}
//: {2}(597,286)(658,286){3}
//: {4}(595,284)(595,249)(606,249){5}
input [15:0] B;    //: /sn:0 {0}(89,381)(128,381){1}
input [15:0] A;    //: /sn:0 {0}(84,200)(130,200){1}
output [15:0] R;    //: /sn:0 {0}(376,288)(421,288){1}
//: {2}(425,288)(464,288){3}
//: {4}(423,286)(423,153)(661,153){5}
output n;    //: /sn:0 /dp:3 {0}(470,213)(541,213){1}
//: {2}(543,211)(543,206)(592,206){3}
//: {4}(596,206)(659,206){5}
//: {6}(594,208)(594,244)(606,244){7}
//: {8}(543,215)(543,249)(551,249){9}
wire w45;    //: /sn:0 {0}(134,346)(214,346){1}
wire w7;    //: /sn:0 {0}(136,175)(213,175){1}
wire w46;    //: /sn:0 {0}(134,336)(214,336){1}
wire w56;    //: /sn:0 {0}(213,255)(136,255){1}
wire w14;    //: /sn:0 {0}(136,225)(213,225){1}
wire w16;    //: /sn:0 {0}(136,205)(213,205){1}
wire w19;    //: /sn:0 {0}(551,314)(535,314)(535,343)(470,343){1}
wire w15;    //: /sn:0 {0}(136,215)(213,215){1}
wire w4;    //: /sn:0 {0}(470,363)(543,363)(543,324)(551,324){1}
wire w38;    //: /sn:0 {0}(134,416)(214,416){1}
wire [15:0] w0;    //: /sn:0 {0}(219,200)(308,200)(308,285)(355,285){1}
wire w3;    //: /sn:0 {0}(136,125)(213,125){1}
wire w37;    //: /sn:0 {0}(134,426)(214,426){1}
wire w34;    //: /sn:0 {0}(136,135)(213,135){1}
wire w43;    //: /sn:0 {0}(134,366)(214,366){1}
wire w21;    //: /sn:0 {0}(470,323)(524,323)(524,304)(551,304){1}
wire [15:0] w58;    //: /sn:0 {0}(220,381)(308,381)(308,290)(355,290){1}
wire w31;    //: /sn:0 {0}(470,223)(540,223)(540,254)(551,254){1}
wire w28;    //: /sn:0 {0}(470,253)(530,253)(530,269)(551,269){1}
wire w36;    //: /sn:0 {0}(134,446)(214,446){1}
wire w41;    //: /sn:0 {0}(134,386)(214,386){1}
wire w20;    //: /sn:0 {0}(470,333)(529,333)(529,309)(551,309){1}
wire w23;    //: /sn:0 {0}(470,303)(516,303)(516,294)(551,294){1}
wire w24;    //: /sn:0 {0}(470,293)(510,293)(510,289)(551,289){1}
wire w1;    //: /sn:0 {0}(136,275)(172,275)(213,275){1}
wire w25;    //: /sn:0 {0}(136,185)(213,185){1}
wire w40;    //: /sn:0 {0}(134,396)(214,396){1}
wire w18;    //: /sn:0 {0}(470,353)(540,353)(540,319)(551,319){1}
wire w8;    //: /sn:0 {0}(136,165)(213,165){1}
wire w30;    //: /sn:0 {0}(470,233)(537,233)(537,259)(551,259){1}
wire w22;    //: /sn:0 {0}(470,313)(520,313)(520,299)(551,299){1}
wire w17;    //: /sn:0 {0}(136,195)(213,195){1}
wire w2;    //: /sn:0 {0}(134,456)(214,456){1}
wire w57;    //: /sn:0 {0}(214,436)(134,436){1}
wire w44;    //: /sn:0 {0}(134,356)(214,356){1}
wire w12;    //: /sn:0 {0}(136,245)(213,245){1}
wire w10;    //: /sn:0 {0}(136,155)(213,155){1}
wire w27;    //: /sn:0 {0}(470,263)(527,263)(527,274)(551,274){1}
wire w13;    //: /sn:0 {0}(136,235)(213,235){1}
wire w48;    //: /sn:0 {0}(134,316)(214,316){1}
wire w5;    //: /sn:0 {0}(136,265)(213,265){1}
wire w33;    //: /sn:0 {0}(136,145)(213,145){1}
wire w47;    //: /sn:0 {0}(134,326)(214,326){1}
wire w29;    //: /sn:0 {0}(470,243)(533,243)(533,264)(551,264){1}
wire w42;    //: /sn:0 {0}(134,376)(214,376){1}
wire w50;    //: /sn:0 {0}(134,306)(214,306){1}
wire w9;    //: /sn:0 {0}(551,284)(510,284)(510,283)(470,283){1}
wire w39;    //: /sn:0 {0}(134,406)(214,406){1}
wire w26;    //: /sn:0 {0}(470,273)(523,273)(523,279)(551,279){1}
//: enddecls

  nor g4 (.I0(n), .I1(z), .Z(p));   //: @(617,247) /sn:0 /w:[ 7 5 0 ]
  //: output g8 (n) @(656,206) /sn:0 /w:[ 5 ]
  //: output g13 (p) @(656,247) /sn:0 /w:[ 1 ]
  //: output g3 (R) @(658,153) /sn:0 /w:[ 5 ]
  //: joint g2 (R) @(423, 288) /w:[ 2 4 1 -1 ]
  or g1 (.I0(w0), .I1(w58), .Z(R));   //: @(366,288) /sn:0 /w:[ 1 1 0 ]
  concat g16 (.I0(w2), .I1(w36), .I2(w57), .I3(w37), .I4(w38), .I5(w39), .I6(w40), .I7(w41), .I8(w42), .I9(w43), .I10(w44), .I11(w45), .I12(w46), .I13(w47), .I14(w48), .I15(w50), .Z(B));   //: @(129,381) /sn:0 /R:2 /w:[ 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:1
  concat g11 (.I0(w4), .I1(w18), .I2(w19), .I3(w20), .I4(w21), .I5(w22), .I6(w23), .I7(w24), .I8(w9), .I9(w26), .I10(w27), .I11(w28), .I12(w29), .I13(w30), .I14(w31), .I15(n), .Z(R));   //: @(465,288) /sn:0 /R:2 /w:[ 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 3 ] /dr:1
  //: joint g6 (n) @(594, 206) /w:[ 4 -1 3 6 ]
  //: joint g9 (z) @(595, 286) /w:[ 2 4 1 -1 ]
  //: input g7 (B) @(87,381) /sn:0 /w:[ 0 ]
  concat g15 (.I0(w1), .I1(w5), .I2(w56), .I3(w12), .I4(w13), .I5(w14), .I6(w15), .I7(w16), .I8(w17), .I9(w25), .I10(w7), .I11(w8), .I12(w10), .I13(w33), .I14(w34), .I15(w3), .Z(A));   //: @(131,200) /sn:0 /R:2 /w:[ 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:1
  concat g17 (.I0(w1), .I1(w5), .I2(w56), .I3(w12), .I4(w13), .I5(w14), .I6(w15), .I7(w16), .I8(w17), .I9(w25), .I10(w7), .I11(w8), .I12(w10), .I13(w33), .I14(w34), .I15(w3), .Z(w0));   //: @(218,200) /sn:0 /w:[ 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 ] /dr:0
  nor g5 (.I0(n), .I1(w31), .I2(w30), .I3(w29), .I4(w28), .I5(w27), .I6(w26), .I7(w9), .I8(w24), .I9(w23), .I10(w22), .I11(w21), .I12(w20), .I13(w19), .I14(w18), .I15(w4), .Z(z));   //: @(562,286) /sn:0 /w:[ 9 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 ]
  //: joint g0 (n) @(543, 213) /w:[ -1 2 1 8 ]
  //: input g22 (A) @(82,200) /sn:0 /w:[ 0 ]
  concat g26 (.I0(w2), .I1(w36), .I2(w57), .I3(w37), .I4(w38), .I5(w39), .I6(w40), .I7(w41), .I8(w42), .I9(w43), .I10(w44), .I11(w45), .I12(w46), .I13(w47), .I14(w48), .I15(w50), .Z(w58));   //: @(219,381) /sn:0 /w:[ 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 ] /dr:0
  //: output g12 (z) @(655,286) /sn:0 /w:[ 3 ]

endmodule

module Soma(B, A, Cin, n, R, o, z, p);
//: interface  /sz:(40, 40) /bd:[ ]
output p;    //: /sn:0 {0}(932,583)(903,583){1}
output z;    //: /sn:0 {0}(931,622)(862,622){1}
//: {2}(860,620)(860,585)(882,585){3}
//: {4}(858,622)(831,622){5}
input [15:0] B;    //: /sn:0 /dp:1 {0}(433,-147)(433,-202){1}
input [15:0] A;    //: /sn:0 {0}(1004,-169)(1004,-194){1}
output [15:0] R;    //: /sn:0 {0}(810,622)(756,622){1}
//: {2}(754,620)(754,576){3}
//: {4}(754,624)(754,676){5}
output o;    //: /sn:0 /dp:1 {0}(934,642)(-77,642)(-77,209)(7,209){1}
input Cin;    //: /sn:0 /dp:3 {0}(1354,195)(1389,195){1}
//: {2}(1393,195)(1407,195){3}
//: {4}(1391,197)(1391,293)(1367,293){5}
output n;    //: /sn:0 {0}(933,546)(862,546){1}
//: {2}(858,546)(831,546){3}
//: {4}(827,546)(218,546)(218,232){5}
//: {6}(829,548)(829,570){7}
//: {8}(860,548)(860,580)(882,580){9}
wire w6;    //: /sn:0 /dp:1 {0}(1178,172)(1178,-115)(488,-115)(488,-141){1}
wire w32;    //: /sn:0 {0}(443,231)(443,267){1}
wire w7;    //: /sn:0 /dp:1 {0}(836,173)(836,116)(948,116)(948,-73)(448,-73)(448,-141){1}
wire c6;    //: /sn:0 {0}(1044,315)(1044,343)(1029,343)(1029,196)(1012,196){1}
wire w16;    //: /sn:0 {0}(1019,-163)(1019,120)(941,120)(941,138)(847,138)(847,173){1}
wire a2;    //: /sn:0 {0}(1189,172)(1189,-144)(1059,-144)(1059,-163){1}
wire p6;    //: /sn:0 {0}(802,267)(802,231){1}
wire Ps;    //: /sn:0 {0}(183,315)(183,347)(161,347)(161,336){1}
wire w4;    //: /sn:0 {0}(699,570)(699,379)(1306,379)(1306,230){1}
wire w15;    //: /sn:0 {0}(1029,-163)(1029,132)(951,132)(951,168)(913,168)(913,173){1}
wire b2;    //: /sn:0 {0}(1255,172)(1255,-148)(1069,-148)(1069,-163){1}
wire w38;    //: /sn:0 /dp:1 {0}(639,231)(639,452)(759,452)(759,570){1}
wire w51;    //: /sn:0 {0}(408,-141)(408,162)(477,162)(477,173){1}
wire w69;    //: /sn:0 {0}(1114,267)(1114,230){1}
wire a4;    //: /sn:0 {0}(488,173)(488,137)(585,137)(585,-7)(979,-7)(979,-163){1}
wire a7;    //: /sn:0 {0}(232,174)(232,-20)(959,-20)(959,-163){1}
wire b11;    //: /sn:0 /dp:1 {0}(554,173)(554,158)(594,158)(594,2)(989,2)(989,-163){1}
wire w0;    //: /sn:0 {0}(-42,118)(-42,192)(7,192){1}
wire w3;    //: /sn:0 {0}(-35,259)(-35,289)(1,289){1}
wire w66;    //: /sn:0 /dp:1 {0}(269,232)(269,504)(799,504)(799,570){1}
wire w64;    //: /sn:0 /dp:1 {0}(53,174)(53,-44)(929,-44)(929,-163){1}
wire w34;    //: /sn:0 /dp:1 {0}(588,231)(588,483)(789,483)(789,570){1}
wire w63;    //: /sn:0 /dp:1 {0}(423,173)(423,133)(575,133)(575,-15)(969,-15)(969,-163){1}
wire w54;    //: /sn:0 {0}(378,-141)(378,-64)(172,-64)(172,174){1}
wire b3;    //: /sn:0 {0}(1243,172)(1243,-122)(498,-122)(498,-141){1}
wire w58;    //: /sn:0 /dp:1 {0}(235,232)(235,530)(819,530)(819,570){1}
wire w28;    //: /sn:0 {0}(739,570)(739,427)(964,427)(964,231){1}
wire w23;    //: /sn:0 {0}(999,-163)(999,11)(602,11)(602,173){1}
wire b6;    //: /sn:0 {0}(901,173)(901,108)(963,108)(963,-82)(458,-82)(458,-141){1}
wire w20;    //: /sn:0 {0}(1340,230)(1340,357)(679,357)(679,570){1}
wire w36;    //: /sn:0 /dp:1 {0}(622,231)(622,461)(769,461)(769,570){1}
wire w1;    //: /sn:0 {0}(710,186)(710,199)(736,199){1}
wire Gs;    //: /sn:0 {0}(142,315)(142,348)(120,348)(120,337){1}
wire b15;    //: /sn:0 /dp:1 {0}(184,174)(184,-28)(949,-28)(949,-163){1}
wire a1;    //: /sn:0 {0}(961,173)(961,142)(1039,142)(1039,-163){1}
wire w65;    //: /sn:0 /dp:1 {0}(252,232)(252,516)(809,516)(809,570){1}
wire a6;    //: /sn:0 {0}(118,174)(118,-38)(939,-38)(939,-163){1}
wire w8;    //: /sn:0 {0}(709,570)(709,391)(1289,391)(1289,230){1}
wire b1;    //: /sn:0 {0}(1290,172)(1290,-128)(508,-128)(508,-141){1}
wire w35;    //: /sn:0 /dp:1 {0}(605,231)(605,471)(779,471)(779,570){1}
wire w40;    //: /sn:0 {0}(43,232)(43,267){1}
wire w30;    //: /sn:0 {0}(749,570)(749,439)(947,439)(947,231){1}
wire w22;    //: /sn:0 {0}(1009,-163)(1009,109)(930,109)(930,137)(782,137)(782,173){1}
wire a0;    //: /sn:0 {0}(1303,172)(1303,-153)(1079,-153)(1079,-163){1}
wire b4;    //: /sn:0 {0}(1099,172)(1099,-108)(478,-108)(478,-141){1}
wire w59;    //: /sn:0 /dp:1 {0}(1124,172)(1124,-139)(1049,-139)(1049,-163){1}
wire b16;    //: /sn:0 {0}(219,174)(219,-58)(388,-58)(388,-141){1}
wire w2;    //: /sn:0 {0}(689,570)(689,368)(1323,368)(1323,230){1}
wire w49;    //: /sn:0 {0}(428,-141)(428,144)(589,144)(589,173){1}
wire cin2;    //: /sn:0 {0}(283,197)(302,197)(302,327)(316,327)(316,315){1}
wire w11;    //: /sn:0 {0}(350,169)(350,189)(377,189){1}
wire w12;    //: /sn:0 {0}(1056,181)(1056,198)(1078,198){1}
wire b8;    //: /sn:0 {0}(948,173)(948,100)(975,100)(975,-93)(468,-93)(468,-141){1}
wire w10;    //: /sn:0 {0}(719,570)(719,404)(998,404)(998,231){1}
wire w13;    //: /sn:0 {0}(729,570)(729,416)(981,416)(981,231){1}
wire w52;    //: /sn:0 {0}(398,-141)(398,173){1}
wire w5;    //: /sn:0 /dp:1 {0}(772,267)(772,231){1}
wire p7;    //: /sn:0 {0}(1144,267)(1144,230){1}
wire w29;    //: /sn:0 {0}(413,231)(413,267){1}
wire p4;    //: /sn:0 {0}(73,267)(73,232){1}
wire w50;    //: /sn:0 {0}(418,-141)(418,156)(542,156)(542,173){1}
wire w9;    //: /sn:0 /dp:1 {0}(107,174)(107,-51)(368,-51)(368,-141){1}
wire b5;    //: /sn:0 {0}(757,173)(757,-64)(438,-64)(438,-141){1}
wire c5;    //: /sn:0 {0}(679,315)(679,325)(666,325)(666,196)(653,196){1}
wire b13;    //: /sn:0 {0}(28,174)(28,-76)(358,-76)(358,-141){1}
//: enddecls

  concat g4 (.I0(a0), .I1(b2), .I2(a2), .I3(w59), .I4(a1), .I5(w15), .I6(w16), .I7(w22), .I8(w23), .I9(b11), .I10(a4), .I11(w63), .I12(a7), .I13(b15), .I14(a6), .I15(w64), .Z(A));   //: @(1004,-168) /sn:0 /R:1 /w:[ 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 ] /dr:0
  led g8 (.I(w0));   //: @(-42,111) /sn:0 /w:[ 0 ] /type:0
  //: input g3 (B) @(433,-204) /sn:0 /R:3 /w:[ 1 ]
  led g13 (.I(w12));   //: @(1056,174) /sn:0 /w:[ 0 ] /type:0
  //: input g2 (A) @(1004,-196) /sn:0 /R:3 /w:[ 1 ]
  //: input g1 (Cin) @(1409,195) /sn:0 /R:2 /w:[ 3 ]
  //: output g16 (n) @(930,546) /sn:0 /w:[ 0 ]
  led g11 (.I(w11));   //: @(350,162) /sn:0 /w:[ 0 ] /type:0
  //: joint g28 (z) @(860, 622) /w:[ 1 2 4 -1 ]
  Somador_CLA_4Bits g10 (.G3(b4), .G2(w6), .G1(b3), .P2(a2), .P3(w59), .P1(b2), .G0(b1), .P0(a0), .Cin(Cin), .C3(w12), .Gs(w69), .Ps(p7), .S3(w8), .S2(w4), .S1(w2), .S0(w20));   //: @(1079, 173) /sz:(274, 56) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Bo2<1 Bo3<1 Bo4<1 Bo5<0 ]
  //: joint g27 (n) @(860, 546) /w:[ 1 -1 2 8 ]
  Somador_CLA_4Bits g19 (.G3(b13), .G2(w9), .G1(w54), .P2(a6), .P3(w64), .P1(b15), .G0(b16), .P0(a7), .Cin(cin2), .O(o), .C3(w0), .Gs(w40), .Ps(p4), .S3(n), .S2(w58), .S1(w65), .S0(w66));   //: @(8, 175) /sz:(274, 56) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>0 Lo0<1 Lo1<1 Bo0<0 Bo1<1 Bo2<5 Bo3<0 Bo4<0 Bo5<0 ]
  concat g6 (.I0(w20), .I1(w2), .I2(w4), .I3(w8), .I4(w10), .I5(w13), .I6(w28), .I7(w30), .I8(w38), .I9(w36), .I10(w35), .I11(w34), .I12(w66), .I13(w65), .I14(w58), .I15(n), .Z(R));   //: @(754,575) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 7 3 ] /dr:0
  //: output g7 (R) @(754,673) /sn:0 /R:3 /w:[ 5 ]
  led g9 (.I(w3));   //: @(-35,252) /sn:0 /w:[ 0 ] /type:0
  //: joint g20 (R) @(754, 622) /w:[ 1 2 -1 4 ]
  //: joint g15 (n) @(829, 546) /w:[ 3 -1 4 6 ]
  //: output g29 (o) @(931,642) /sn:0 /w:[ 0 ]
  nor g25 (.I0(n), .I1(z), .Z(p));   //: @(893,583) /sn:0 /w:[ 9 3 1 ]
  Somador_CLA_4Bits g17 (.G3(b5), .G2(w7), .G1(b6), .P2(w16), .P3(w22), .P1(w15), .G0(b8), .P0(a1), .Cin(c6), .C3(w1), .Gs(w5), .Ps(p6), .S3(w30), .S2(w28), .S1(w13), .S0(w10));   //: @(737, 174) /sz:(274, 56) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>1 Ti4>1 Ti5>1 Ti6>0 Ti7>0 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Bo2<1 Bo3<1 Bo4<1 Bo5<1 ]
  concat g5 (.I0(b1), .I1(b3), .I2(w6), .I3(b4), .I4(b8), .I5(b6), .I6(w7), .I7(b5), .I8(w49), .I9(w50), .I10(w51), .I11(w52), .I12(b16), .I13(w54), .I14(w9), .I15(b13), .Z(B));   //: @(433,-146) /sn:0 /R:1 /w:[ 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 ] /dr:0
  //: output g24 (z) @(928,622) /sn:0 /w:[ 0 ]
  led g21 (.I(Ps));   //: @(161,329) /sn:0 /w:[ 1 ] /type:0
  nor g23 (.I0(R), .Z(z));   //: @(821,622) /sn:0 /w:[ 0 5 ]
  //: output g26 (p) @(929,583) /sn:0 /w:[ 0 ]
  //: joint g0 (Cin) @(1391, 195) /w:[ 2 -1 1 4 ]
  led g22 (.I(Gs));   //: @(120,330) /sn:0 /w:[ 1 ] /type:0
  Somador_CLA_4Bits g18 (.G3(w52), .G2(w51), .G1(w50), .P2(a4), .P3(w63), .P1(b11), .G0(w49), .P0(w23), .Cin(c5), .C3(w11), .Gs(w29), .Ps(w32), .S3(w34), .S2(w35), .S1(w36), .S0(w38));   //: @(378, 174) /sz:(274, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>0 Ti4>0 Ti5>0 Ti6>1 Ti7>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Bo2<0 Bo3<0 Bo4<0 Bo5<0 ]
  led g12 (.I(w1));   //: @(710,179) /sn:0 /w:[ 0 ] /type:0
  CLA g91 (.G3(w40), .P3(p4), .G2(w29), .P2(w32), .G1(w5), .P1(p6), .G0(w69), .P0(p7), .Cin(Cin), .C3(w3), .Ps(Ps), .Gs(Gs), .C2(cin2), .C1(c5), .C0(c6));   //: @(2, 268) /sz:(1364, 46) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>1 Ti3>1 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>5 Lo0<1 Bo0<0 Bo1<0 Bo2<1 Bo3<0 Bo4<0 ]

endmodule

module SUB(B, A, Cin, n, R, o, z, p);
//: interface  /sz:(40, 40) /bd:[ ]
output p;    //: /sn:0 {0}(546,459)(517,459){1}
input [15:0] B;    //: /sn:0 /dp:1 {0}(47,-329)(47,-351){1}
output z;    //: /sn:0 {0}(545,498)(476,498){1}
//: {2}(474,496)(474,461)(496,461){3}
//: {4}(472,498)(445,498){5}
input [15:0] A;    //: /sn:0 {0}(618,-293)(618,-344){1}
output [15:0] R;    //: /sn:0 {0}(424,498)(370,498){1}
//: {2}(368,496)(368,452){3}
//: {4}(368,500)(368,552){5}
output o;    //: /sn:0 {0}(548,518)(-463,518)(-463,85)(-379,85){1}
input Cin;    //: /sn:0 {0}(968,71)(1003,71){1}
//: {2}(1007,71)(1021,71){3}
//: {4}(1005,73)(1005,169)(981,169){5}
output n;    //: /sn:0 {0}(547,422)(476,422){1}
//: {2}(472,422)(445,422){3}
//: {4}(441,422)(-168,422)(-168,108){5}
//: {6}(443,424)(443,446){7}
//: {8}(474,424)(474,456)(496,456){9}
wire w32;    //: /sn:0 {0}(57,107)(57,143){1}
wire w6;    //: /sn:0 {0}(792,48)(792,-239)(102,-239)(102,-265){1}
wire w7;    //: /sn:0 {0}(450,49)(450,-8)(562,-8)(562,-197)(62,-197)(62,-265){1}
wire c6;    //: /sn:0 {0}(658,191)(658,219)(643,219)(643,72)(626,72){1}
wire Ps;    //: /sn:0 {0}(-203,191)(-203,223)(-225,223)(-225,212){1}
wire p6;    //: /sn:0 {0}(416,143)(416,107){1}
wire w16;    //: /sn:0 {0}(633,-287)(633,-4)(555,-4)(555,14)(461,14)(461,49){1}
wire a2;    //: /sn:0 {0}(803,48)(803,-268)(673,-268)(673,-287){1}
wire w4;    //: /sn:0 {0}(313,446)(313,255)(920,255)(920,106){1}
wire w15;    //: /sn:0 {0}(643,-287)(643,8)(565,8)(565,44)(527,44)(527,49){1}
wire b2;    //: /sn:0 {0}(869,48)(869,-272)(683,-272)(683,-287){1}
wire w38;    //: /sn:0 {0}(253,107)(253,328)(373,328)(373,446){1}
wire w51;    //: /sn:0 {0}(22,-265)(22,38)(91,38)(91,49){1}
wire w69;    //: /sn:0 {0}(728,143)(728,106){1}
wire a7;    //: /sn:0 {0}(-154,50)(-154,-144)(573,-144)(573,-287){1}
wire a4;    //: /sn:0 {0}(102,49)(102,13)(199,13)(199,-131)(593,-131)(593,-287){1}
wire w3;    //: /sn:0 {0}(-421,135)(-421,165)(-385,165){1}
wire b11;    //: /sn:0 {0}(168,49)(168,34)(208,34)(208,-122)(603,-122)(603,-287){1}
wire w0;    //: /sn:0 {0}(-428,-6)(-428,68)(-379,68){1}
wire w66;    //: /sn:0 {0}(-117,108)(-117,380)(413,380)(413,446){1}
wire w64;    //: /sn:0 {0}(-333,50)(-333,-168)(543,-168)(543,-287){1}
wire w34;    //: /sn:0 {0}(202,107)(202,359)(403,359)(403,446){1}
wire w63;    //: /sn:0 {0}(37,49)(37,9)(189,9)(189,-139)(583,-139)(583,-287){1}
wire w54;    //: /sn:0 {0}(-8,-265)(-8,-188)(-214,-188)(-214,50){1}
wire b3;    //: /sn:0 {0}(857,48)(857,-246)(112,-246)(112,-265){1}
wire w58;    //: /sn:0 {0}(-151,108)(-151,406)(433,406)(433,446){1}
wire w28;    //: /sn:0 {0}(353,446)(353,303)(578,303)(578,107){1}
wire b6;    //: /sn:0 {0}(515,49)(515,-16)(577,-16)(577,-206)(72,-206)(72,-265){1}
wire w36;    //: /sn:0 {0}(236,107)(236,337)(383,337)(383,446){1}
wire w20;    //: /sn:0 {0}(954,106)(954,233)(293,233)(293,446){1}
wire w23;    //: /sn:0 {0}(613,-287)(613,-113)(216,-113)(216,49){1}
wire w1;    //: /sn:0 {0}(324,62)(324,75)(350,75){1}
wire Gs;    //: /sn:0 {0}(-244,191)(-244,224)(-266,224)(-266,213){1}
wire b15;    //: /sn:0 {0}(-202,50)(-202,-152)(563,-152)(563,-287){1}
wire w65;    //: /sn:0 {0}(-134,108)(-134,392)(423,392)(423,446){1}
wire a6;    //: /sn:0 {0}(-268,50)(-268,-162)(553,-162)(553,-287){1}
wire a1;    //: /sn:0 {0}(575,49)(575,18)(653,18)(653,-287){1}
wire [15:0] w18;    //: /sn:0 /dp:1 {0}(47,-313)(47,-271){1}
wire w35;    //: /sn:0 {0}(219,107)(219,347)(393,347)(393,446){1}
wire w40;    //: /sn:0 {0}(-343,108)(-343,143){1}
wire w8;    //: /sn:0 {0}(323,446)(323,267)(903,267)(903,106){1}
wire b1;    //: /sn:0 {0}(904,48)(904,-252)(122,-252)(122,-265){1}
wire w30;    //: /sn:0 {0}(363,446)(363,315)(561,315)(561,107){1}
wire b4;    //: /sn:0 {0}(713,48)(713,-232)(92,-232)(92,-265){1}
wire w22;    //: /sn:0 {0}(623,-287)(623,-15)(544,-15)(544,13)(396,13)(396,49){1}
wire a0;    //: /sn:0 {0}(917,48)(917,-277)(693,-277)(693,-287){1}
wire w59;    //: /sn:0 {0}(738,48)(738,-263)(663,-263)(663,-287){1}
wire b16;    //: /sn:0 {0}(-167,50)(-167,-182)(2,-182)(2,-265){1}
wire w49;    //: /sn:0 {0}(42,-265)(42,20)(203,20)(203,49){1}
wire cin2;    //: /sn:0 {0}(-103,73)(-84,73)(-84,203)(-70,203)(-70,191){1}
wire w2;    //: /sn:0 {0}(303,446)(303,244)(937,244)(937,106){1}
wire w11;    //: /sn:0 {0}(-36,45)(-36,65)(-9,65){1}
wire w12;    //: /sn:0 {0}(670,57)(670,74)(692,74){1}
wire b8;    //: /sn:0 {0}(562,49)(562,-24)(589,-24)(589,-217)(82,-217)(82,-265){1}
wire w10;    //: /sn:0 {0}(333,446)(333,280)(612,280)(612,107){1}
wire w13;    //: /sn:0 {0}(343,446)(343,292)(595,292)(595,107){1}
wire w52;    //: /sn:0 {0}(12,-265)(12,49){1}
wire w5;    //: /sn:0 {0}(386,143)(386,107){1}
wire p7;    //: /sn:0 {0}(758,143)(758,106){1}
wire w29;    //: /sn:0 {0}(27,107)(27,143){1}
wire p4;    //: /sn:0 {0}(-313,143)(-313,108){1}
wire w50;    //: /sn:0 {0}(32,-265)(32,32)(156,32)(156,49){1}
wire w9;    //: /sn:0 {0}(-279,50)(-279,-175)(-18,-175)(-18,-265){1}
wire c5;    //: /sn:0 {0}(293,191)(293,201)(280,201)(280,72)(267,72){1}
wire b5;    //: /sn:0 {0}(371,49)(371,-188)(52,-188)(52,-265){1}
wire b13;    //: /sn:0 {0}(-358,50)(-358,-200)(-28,-200)(-28,-265){1}
//: enddecls

  concat g4 (.I0(a0), .I1(b2), .I2(a2), .I3(w59), .I4(a1), .I5(w15), .I6(w16), .I7(w22), .I8(w23), .I9(b11), .I10(a4), .I11(w63), .I12(a7), .I13(b15), .I14(a6), .I15(w64), .Z(A));   //: @(618,-292) /sn:0 /R:1 /w:[ 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 ] /dr:0
  led g8 (.I(w0));   //: @(-428,-13) /sn:0 /w:[ 0 ] /type:0
  //: input g3 (B) @(47,-353) /sn:0 /R:3 /w:[ 1 ]
  led g13 (.I(w12));   //: @(670,50) /sn:0 /w:[ 0 ] /type:0
  //: input g2 (A) @(618,-346) /sn:0 /R:3 /w:[ 1 ]
  //: input g1 (Cin) @(1023,71) /sn:0 /R:2 /w:[ 3 ]
  //: output g16 (n) @(544,422) /sn:0 /w:[ 0 ]
  led g11 (.I(w11));   //: @(-36,38) /sn:0 /w:[ 0 ] /type:0
  //: joint g28 (z) @(474, 498) /w:[ 1 2 4 -1 ]
  Somador_CLA_4Bits g10 (.G3(b4), .G2(w6), .G1(b3), .P2(a2), .P3(w59), .P1(b2), .G0(b1), .P0(a0), .Cin(Cin), .C3(w12), .Gs(w69), .Ps(p7), .S3(w8), .S2(w4), .S1(w2), .S0(w20));   //: @(693, 49) /sz:(274, 56) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Bo2<1 Bo3<1 Bo4<1 Bo5<0 ]
  //: joint g27 (n) @(474, 422) /w:[ 1 -1 2 8 ]
  Somador_CLA_4Bits g19 (.G3(b13), .G2(w9), .G1(w54), .P2(a6), .P3(w64), .P1(b15), .G0(b16), .P0(a7), .Cin(cin2), .O(o), .C3(w0), .Gs(w40), .Ps(p4), .S3(n), .S2(w58), .S1(w65), .S0(w66));   //: @(-378, 51) /sz:(274, 56) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>0 Lo0<1 Lo1<1 Bo0<0 Bo1<1 Bo2<5 Bo3<0 Bo4<0 Bo5<0 ]
  concat g6 (.I0(w20), .I1(w2), .I2(w4), .I3(w8), .I4(w10), .I5(w13), .I6(w28), .I7(w30), .I8(w38), .I9(w36), .I10(w35), .I11(w34), .I12(w66), .I13(w65), .I14(w58), .I15(n), .Z(R));   //: @(368,451) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 7 3 ] /dr:0
  //: output g7 (R) @(368,549) /sn:0 /R:3 /w:[ 5 ]
  led g9 (.I(w3));   //: @(-421,128) /sn:0 /w:[ 0 ] /type:0
  //: joint g20 (R) @(368, 498) /w:[ 1 2 -1 4 ]
  //: joint g15 (n) @(443, 422) /w:[ 3 -1 4 6 ]
  //: output g29 (o) @(545,518) /sn:0 /w:[ 0 ]
  nor g25 (.I0(n), .I1(z), .Z(p));   //: @(507,459) /sn:0 /w:[ 9 3 1 ]
  Somador_CLA_4Bits g17 (.G3(b5), .G2(w7), .G1(b6), .P2(w16), .P3(w22), .P1(w15), .G0(b8), .P0(a1), .Cin(c6), .C3(w1), .Gs(w5), .Ps(p6), .S3(w30), .S2(w28), .S1(w13), .S0(w10));   //: @(351, 50) /sz:(274, 56) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>1 Ti4>1 Ti5>1 Ti6>0 Ti7>0 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Bo2<1 Bo3<1 Bo4<1 Bo5<1 ]
  not g14 (.I(B), .Z(w18));   //: @(47,-323) /sn:0 /R:3 /w:[ 0 0 ]
  concat g5 (.I0(b1), .I1(b3), .I2(w6), .I3(b4), .I4(b8), .I5(b6), .I6(w7), .I7(b5), .I8(w49), .I9(w50), .I10(w51), .I11(w52), .I12(b16), .I13(w54), .I14(w9), .I15(b13), .Z(w18));   //: @(47,-270) /sn:0 /R:1 /w:[ 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1 1 1 ] /dr:0
  //: output g24 (z) @(542,498) /sn:0 /w:[ 0 ]
  led g21 (.I(Ps));   //: @(-225,205) /sn:0 /w:[ 1 ] /type:0
  nor g23 (.I0(R), .Z(z));   //: @(435,498) /sn:0 /w:[ 0 5 ]
  //: output g26 (p) @(543,459) /sn:0 /w:[ 0 ]
  //: joint g0 (Cin) @(1005, 71) /w:[ 2 -1 1 4 ]
  led g22 (.I(Gs));   //: @(-266,206) /sn:0 /w:[ 1 ] /type:0
  Somador_CLA_4Bits g18 (.G3(w52), .G2(w51), .G1(w50), .P2(a4), .P3(w63), .P1(b11), .G0(w49), .P0(w23), .Cin(c5), .C3(w11), .Gs(w29), .Ps(w32), .S3(w34), .S2(w35), .S1(w36), .S0(w38));   //: @(-8, 50) /sz:(274, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>0 Ti4>0 Ti5>0 Ti6>1 Ti7>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Bo2<0 Bo3<0 Bo4<0 Bo5<0 ]
  led g12 (.I(w1));   //: @(324,55) /sn:0 /w:[ 0 ] /type:0
  CLA g91 (.G3(w40), .P3(p4), .G2(w29), .P2(w32), .G1(w5), .P1(p6), .G0(w69), .P0(p7), .Cin(Cin), .C3(w3), .Ps(Ps), .Gs(Gs), .C2(cin2), .C1(c5), .C0(c6));   //: @(-384, 144) /sz:(1364, 46) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>1 Ti3>1 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>5 Lo0<1 Bo0<0 Bo1<0 Bo2<1 Bo3<0 Bo4<0 ]

endmodule

module REGISTRADORES(RegBusB, DataOutBusB, DataOutBusA, LoadReg, RegDst, CLK, RegBusA, Reset, R);
//: interface  /sz:(40, 40) /bd:[ ]
input LoadReg;    //: /sn:0 {0}(80,199)(90,199)(90,472)(147,472)(147,461){1}
input [3:0] RegBusA;    //: /sn:0 {0}(86,53)(593,53)(593,272)(573,272)(573,262){1}
input [15:0] R;    //: /sn:0 {0}(310,268)(310,261)(251,261){1}
//: {2}(249,259)(249,214){3}
//: {4}(251,212)(309,212)(309,221){5}
//: {6}(249,210)(249,173){7}
//: {8}(251,171)(309,171)(309,178){9}
//: {10}(249,169)(249,119){11}
//: {12}(251,117)(308,117)(308,135){13}
//: {14}(247,117)(83,117){15}
//: {16}(249,263)(249,303){17}
//: {18}(251,305)(312,305)(312,311){19}
//: {20}(249,307)(249,345){21}
//: {22}(251,347)(312,347)(312,352){23}
//: {24}(249,349)(249,386){25}
//: {26}(251,388)(313,388)(313,392){27}
//: {28}(249,390)(249,427){29}
//: {30}(251,429)(313,429)(313,437){31}
//: {32}(249,431)(249,473){33}
//: {34}(251,475)(313,475)(313,483){35}
//: {36}(249,477)(249,520){37}
//: {38}(251,522)(315,522)(315,533){39}
//: {40}(249,524)(249,566){41}
//: {42}(251,568)(316,568)(316,576){43}
//: {44}(249,570)(249,613)(317,613)(317,621){45}
output [15:0] DataOutBusA;    //: /sn:0 {0}(641,239)(586,239){1}
output [15:0] DataOutBusB;    //: /sn:0 /dp:1 {0}(590,361)(648,361){1}
input [3:0] RegDst;    //: /sn:0 {0}(82,172)(100,172)(100,439)(134,439){1}
input CLK;    //: /sn:0 {0}(83,145)(259,145){1}
//: {2}(263,145)(271,145){3}
//: {4}(261,147)(261,186){5}
//: {6}(263,188)(272,188){7}
//: {8}(261,190)(261,229){9}
//: {10}(263,231)(272,231){11}
//: {12}(261,233)(261,276){13}
//: {14}(263,278)(273,278){15}
//: {16}(261,280)(261,319){17}
//: {18}(263,321)(275,321){19}
//: {20}(261,323)(261,360){21}
//: {22}(263,362)(275,362){23}
//: {24}(261,364)(261,400){25}
//: {26}(263,402)(276,402){27}
//: {28}(261,404)(261,445){29}
//: {30}(263,447)(276,447){31}
//: {32}(261,449)(261,491){33}
//: {34}(263,493)(276,493){35}
//: {36}(261,495)(261,541){37}
//: {38}(263,543)(278,543){39}
//: {40}(261,545)(261,584){41}
//: {42}(263,586)(279,586){43}
//: {44}(261,588)(261,631)(280,631){45}
input Reset;    //: /sn:0 {0}(85,97)(373,97)(373,138){1}
//: {2}(371,140)(347,140){3}
//: {4}(373,142)(373,181){5}
//: {6}(371,183)(348,183){7}
//: {8}(373,185)(373,224){9}
//: {10}(371,226)(348,226){11}
//: {12}(373,228)(373,271){13}
//: {14}(371,273)(349,273){15}
//: {16}(373,275)(373,314){17}
//: {18}(371,316)(351,316){19}
//: {20}(373,318)(373,355){21}
//: {22}(371,357)(351,357){23}
//: {24}(373,359)(373,395){25}
//: {26}(371,397)(352,397){27}
//: {28}(373,399)(373,440){29}
//: {30}(371,442)(352,442){31}
//: {32}(373,444)(373,486){33}
//: {34}(371,488)(352,488){35}
//: {36}(373,490)(373,536){37}
//: {38}(371,538)(354,538){39}
//: {40}(373,540)(373,579){41}
//: {42}(371,581)(355,581){43}
//: {44}(373,583)(373,626)(356,626){45}
input [3:0] RegBusB;    //: /sn:0 {0}(85,75)(605,75)(605,394)(577,394)(577,384){1}
wire [15:0] w45;    //: /sn:0 {0}(315,554)(315,560)(461,560)(461,255)(491,255){1}
//: {2}(495,255)(557,255){3}
//: {4}(493,257)(493,377)(561,377){5}
wire [15:0] w73;    //: /sn:0 /dp:1 {0}(557,264)(481,264){1}
//: {2}(477,264)(472,264)(472,653)(317,653)(317,642){3}
//: {4}(479,266)(479,386)(561,386){5}
wire w96;    //: /sn:0 {0}(163,441)(208,441)(208,417)(357,417)(357,407)(352,407){1}
wire w7;    //: /sn:0 /dp:1 {0}(348,193)(355,193)(355,203)(181,203)(181,418)(163,418){1}
wire [15:0] w60;    //: /sn:0 {0}(557,213)(554,213){1}
//: {2}(550,213)(430,213)(430,164)(308,164)(308,156){3}
//: {4}(552,215)(552,335)(561,335){5}
wire w99;    //: /sn:0 {0}(163,455)(189,455)(189,531)(358,531)(358,548)(354,548){1}
wire w16;    //: /sn:0 /dp:1 {0}(348,236)(354,236)(354,247)(188,247)(188,422)(163,422){1}
wire [15:0] w0;    //: /sn:0 {0}(309,242)(309,255)(420,255)(420,222)(537,222){1}
//: {2}(541,222)(557,222){3}
//: {4}(539,224)(539,344)(561,344){5}
wire w97;    //: /sn:0 {0}(163,445)(201,445)(201,464)(358,464)(358,452)(352,452){1}
wire [15:0] w66;    //: /sn:0 {0}(557,241)(515,241){1}
//: {2}(511,241)(445,241)(445,424)(313,424)(313,413){3}
//: {4}(513,243)(513,363)(561,363){5}
wire [15:0] w64;    //: /sn:0 {0}(557,232)(528,232){1}
//: {2}(524,232)(436,232)(436,342)(312,342)(312,332){3}
//: {4}(526,234)(526,354)(561,354){5}
wire w90;    //: /sn:0 {0}(163,413)(176,413)(176,159)(354,159)(354,150)(347,150){1}
wire [15:0] w28;    //: /sn:0 {0}(557,245)(509,245){1}
//: {2}(505,245)(450,245)(450,469)(313,469)(313,458){3}
//: {4}(507,247)(507,367)(561,367){5}
wire [15:0] w65;    //: /sn:0 {0}(557,236)(522,236){1}
//: {2}(518,236)(441,236)(441,381)(312,381)(312,373){3}
//: {4}(520,238)(520,358)(561,358){5}
wire [15:0] w40;    //: /sn:0 {0}(316,597)(316,603)(466,603)(466,259)(484,259){1}
//: {2}(488,259)(557,259){3}
//: {4}(486,261)(486,381)(561,381){5}
wire w101;    //: /sn:0 {0}(163,464)(178,464)(178,617)(366,617)(366,636)(356,636){1}
wire [15:0] w2;    //: /sn:0 /dp:1 {0}(557,227)(535,227){1}
//: {2}(531,227)(430,227)(430,298)(310,298)(310,289){3}
//: {4}(533,229)(533,349)(561,349){5}
wire w12;    //: /sn:0 /dp:1 {0}(349,283)(360,283)(360,294)(192,294)(192,427)(163,427){1}
wire w94;    //: /sn:0 {0}(163,432)(197,432)(197,337)(361,337)(361,326)(351,326){1}
wire [15:0] w5;    //: /sn:0 /dp:1 {0}(309,199)(309,207)(428,207)(428,218)(544,218){1}
//: {2}(548,218)(557,218){3}
//: {4}(546,220)(546,340)(561,340){5}
wire w95;    //: /sn:0 {0}(163,436)(203,436)(203,377)(361,377)(361,367)(351,367){1}
wire w52;    //: /sn:0 /dp:1 {0}(352,498)(359,498)(359,483)(191,483)(191,450)(163,450){1}
wire [15:0] w50;    //: /sn:0 {0}(313,504)(313,515)(454,515)(454,250)(498,250){1}
//: {2}(502,250)(557,250){3}
//: {4}(500,252)(500,372)(561,372){5}
wire w42;    //: /sn:0 /dp:1 {0}(355,591)(362,591)(362,574)(183,574)(183,459)(163,459){1}
//: enddecls

  //: joint g61 (Reset) @(373, 357) /w:[ -1 21 22 24 ]
  register REG2 (.Q(w5), .D(R), .EN(w7), .CLR(Reset), .CK(CLK));   //: @(309,188) /w:[ 0 9 0 7 7 ]
  register REG7 (.Q(w66), .D(R), .EN(w96), .CLR(Reset), .CK(CLK));   //: @(313,402) /w:[ 3 27 1 27 27 ]
  //: joint g58 (Reset) @(373, 488) /w:[ -1 33 34 36 ]
  //: input g55 (RegBusB) @(83,75) /sn:0 /w:[ 0 ]
  //: joint g51 (CLK) @(261, 493) /w:[ 34 33 -1 36 ]
  //: joint g37 (R) @(249, 429) /w:[ 30 29 -1 32 ]
  //: joint g34 (R) @(249, 305) /w:[ 18 17 -1 20 ]
  //: joint g13 (w60) @(552, 213) /w:[ 1 -1 2 4 ]
  //: joint g65 (Reset) @(373, 183) /w:[ -1 5 6 8 ]
  register REG12 (.Q(w73), .D(R), .EN(w101), .CLR(Reset), .CK(CLK));   //: @(317,631) /w:[ 3 45 1 45 45 ]
  //: joint g59 (Reset) @(373, 442) /w:[ -1 29 30 32 ]
  //: joint g64 (Reset) @(373, 226) /w:[ -1 9 10 12 ]
  //: joint g16 (w5) @(546, 218) /w:[ 2 -1 1 4 ]
  //: joint g50 (CLK) @(261, 447) /w:[ 30 29 -1 32 ]
  //: output g28 (DataOutBusB) @(645,361) /sn:0 /w:[ 1 ]
  register REG4 (.Q(w2), .D(R), .EN(w12), .CLR(Reset), .CK(CLK));   //: @(310,278) /w:[ 3 0 0 15 15 ]
  //: joint g32 (R) @(249, 171) /w:[ 8 10 -1 7 ]
  //: output g27 (DataOutBusA) @(638,239) /sn:0 /w:[ 0 ]
  //: joint g19 (w64) @(526, 232) /w:[ 1 -1 2 4 ]
  //: joint g38 (R) @(249, 475) /w:[ 34 33 -1 36 ]
  //: joint g57 (Reset) @(373, 538) /w:[ -1 37 38 40 ]
  //: joint g53 (CLK) @(261, 586) /w:[ 42 41 -1 44 ]
  //: joint g31 (R) @(249, 117) /w:[ 12 -1 14 11 ]
  //: joint g20 (w65) @(520, 236) /w:[ 1 -1 2 4 ]
  mux g15 (.I0(w60), .I1(w5), .I2(w0), .I3(w2), .I4(w64), .I5(w65), .I6(w66), .I7(w28), .I8(w50), .I9(w45), .I10(w40), .I11(w73), .S(RegBusB), .Z(DataOutBusB));   //: @(577,361) /sn:0 /R:1 /w:[ 5 5 5 5 5 5 5 5 5 5 5 5 1 0 ] /ss:0 /do:0
  //: input g68 (LoadReg) @(78,199) /sn:0 /w:[ 0 ]
  //: joint g67 (Reset) @(373, 140) /w:[ -1 1 2 4 ]
  //: joint g39 (R) @(249, 522) /w:[ 38 37 -1 40 ]
  register REG1 (.Q(w60), .D(R), .EN(w90), .CLR(Reset), .CK(CLK));   //: @(308,145) /w:[ 3 13 1 3 3 ]
  register REG9 (.Q(w50), .D(R), .EN(w52), .CLR(Reset), .CK(CLK));   //: @(313,493) /w:[ 0 35 0 35 35 ]
  //: joint g48 (CLK) @(261, 362) /w:[ 22 21 -1 24 ]
  //: joint g43 (CLK) @(261, 145) /w:[ 2 -1 1 4 ]
  register REG8 (.Q(w28), .D(R), .EN(w97), .CLR(Reset), .CK(CLK));   //: @(313,447) /w:[ 3 31 1 31 31 ]
  //: joint g62 (Reset) @(373, 316) /w:[ -1 17 18 20 ]
  //: input g29 (RegDst) @(80,172) /sn:0 /w:[ 0 ]
  //: joint g25 (w40) @(486, 259) /w:[ 2 -1 1 4 ]
  //: joint g17 (w0) @(539, 222) /w:[ 2 -1 1 4 ]
  //: joint g63 (Reset) @(373, 273) /w:[ -1 13 14 16 ]
  //: joint g52 (CLK) @(261, 543) /w:[ 38 37 -1 40 ]
  //: input g42 (CLK) @(81,145) /sn:0 /w:[ 0 ]
  register REG3 (.Q(w0), .D(R), .EN(w16), .CLR(Reset), .CK(CLK));   //: @(309,231) /w:[ 0 5 0 11 11 ]
  register REG5 (.Q(w64), .D(R), .EN(w94), .CLR(Reset), .CK(CLK));   //: @(312,321) /w:[ 3 19 1 19 19 ]
  //: joint g56 (Reset) @(373, 581) /w:[ -1 41 42 44 ]
  demux g14 (.I(RegDst), .E(LoadReg), .Z0(w90), .Z1(w7), .Z2(w16), .Z3(w12), .Z4(w94), .Z5(w95), .Z6(w96), .Z7(w97), .Z8(w52), .Z9(w99), .Z10(w42), .Z11(w101));   //: @(147,439) /sn:0 /R:1 /w:[ 1 1 0 1 1 1 0 0 0 0 1 0 1 0 ]
  //: joint g47 (CLK) @(261, 321) /w:[ 18 17 -1 20 ]
  //: joint g44 (CLK) @(261, 188) /w:[ 6 5 -1 8 ]
  //: joint g36 (R) @(249, 388) /w:[ 26 25 -1 28 ]
  //: joint g24 (w45) @(493, 255) /w:[ 2 -1 1 4 ]
  //: joint g21 (w66) @(513, 241) /w:[ 1 -1 2 4 ]
  //: joint g41 (R) @(249, 261) /w:[ 1 2 -1 16 ]
  //: joint g23 (w50) @(500, 250) /w:[ 2 -1 1 4 ]
  register REG11 (.Q(w40), .D(R), .EN(w42), .CLR(Reset), .CK(CLK));   //: @(316,586) /w:[ 0 43 0 43 43 ]
  //: joint g60 (Reset) @(373, 397) /w:[ -1 25 26 28 ]
  //: input g54 (RegBusA) @(84,53) /sn:0 /w:[ 0 ]
  //: joint g40 (R) @(249, 568) /w:[ 42 41 -1 44 ]
  register REG6 (.Q(w65), .D(R), .EN(w95), .CLR(Reset), .CK(CLK));   //: @(312,362) /w:[ 3 23 1 23 23 ]
  //: joint g46 (CLK) @(261, 278) /w:[ 14 13 -1 16 ]
  //: joint g45 (CLK) @(261, 231) /w:[ 10 9 -1 12 ]
  //: joint g35 (R) @(249, 347) /w:[ 22 21 -1 24 ]
  //: joint g26 (w73) @(479, 264) /w:[ 1 -1 2 4 ]
  //: joint g22 (w28) @(507, 245) /w:[ 1 -1 2 4 ]
  //: input g66 (Reset) @(83,97) /sn:0 /w:[ 0 ]
  //: joint g18 (w2) @(533, 227) /w:[ 1 -1 2 4 ]
  mux g12 (.I0(w60), .I1(w5), .I2(w0), .I3(w2), .I4(w64), .I5(w65), .I6(w66), .I7(w28), .I8(w50), .I9(w45), .I10(w40), .I11(w73), .S(RegBusA), .Z(DataOutBusA));   //: @(573,239) /sn:0 /R:1 /w:[ 0 3 3 0 0 0 0 0 3 3 3 0 1 1 ] /ss:0 /do:0
  //: joint g33 (R) @(249, 212) /w:[ 4 6 -1 3 ]
  //: input g30 (R) @(81,117) /sn:0 /w:[ 15 ]
  register REG10 (.Q(w45), .D(R), .EN(w99), .CLR(Reset), .CK(CLK));   //: @(315,543) /w:[ 0 39 1 39 39 ]
  //: joint g49 (CLK) @(261, 402) /w:[ 26 25 -1 28 ]

endmodule

module REGSTAT(en, z, p, o, CLK, n, S);
//: interface  /sz:(40, 40) /bd:[ ]
output p;    //: /sn:0 {0}(334,294)(334,256){1}
output z;    //: /sn:0 {0}(324,294)(324,256){1}
supply1 w0;    //: /sn:0 {0}(394,156)(394,192)(368,192){1}
input en;    //: /sn:0 {0}(422,202)(368,202){1}
output o;    //: /sn:0 {0}(344,294)(344,256){1}
input CLK;    //: /sn:0 {0}(265,197)(292,197){1}
output n;    //: /sn:0 {0}(314,294)(314,256){1}
input [3:0] S;    //: /sn:0 {0}(261,156)(329,156)(329,187){1}
wire [3:0] sta;    //: /sn:0 {0}(329,250)(329,208){1}
//: enddecls

  //: input g8 (en) @(424,202) /sn:0 /R:2 /w:[ 0 ]
  //: output g4 (z) @(324,291) /sn:0 /R:3 /w:[ 0 ]
  //: output g3 (p) @(334,291) /sn:0 /R:3 /w:[ 0 ]
  //: output g2 (o) @(344,291) /sn:0 /R:3 /w:[ 0 ]
  concat g1 (.I0(o), .I1(p), .I2(z), .I3(n), .Z(sta));   //: @(329,251) /sn:0 /R:1 /w:[ 1 1 1 1 0 ] /dr:0
  register REGSTAT (.Q(sta), .D(S), .EN(en), .CLR(w0), .CK(CLK));   //: @(329,197) /w:[ 1 1 1 1 1 ]
  //: input g9 (CLK) @(263,197) /sn:0 /w:[ 0 ]
  //: supply1 g7 (w0) @(405,156) /sn:0 /w:[ 0 ]
  //: output g5 (n) @(314,291) /sn:0 /R:3 /w:[ 0 ]
  //: input g0 (S) @(259,156) /sn:0 /w:[ 0 ]

endmodule

module Somador_CLA_4Bits(P2, S2, G3, S1, S0, Ps, G1, G0, P0, P3, P1, Cin, O, C3, S3, Gs, G2);
//: interface  /sz:(40, 40) /bd:[ ]
output S1;    //: /sn:0 {0}(577,447)(577,312){1}
input G2;    //: /sn:0 {0}(320,91)(320,202){1}
//: {2}(322,204)(337,204)(337,218){3}
//: {4}(320,206)(320,216){5}
output Ps;    //: /sn:0 {0}(206,441)(206,407){1}
input P1;    //: /sn:0 {0}(535,90)(535,199){1}
//: {2}(533,201)(507,201)(507,219){3}
//: {4}(535,203)(535,220){5}
output C3;    //: /sn:0 /dp:1 {0}(79,381)(99,381){1}
//: {2}(103,381)(126,381){3}
//: {4}(101,379)(101,302){5}
input G0;    //: /sn:0 {0}(659,90)(659,203){1}
//: {2}(661,205)(680,205)(680,217){3}
//: {4}(659,207)(659,217){5}
output Gs;    //: /sn:0 {0}(188,442)(188,407){1}
output S0;    //: /sn:0 /dp:1 {0}(709,324)(709,343)(696,343)(696,447){1}
input P3;    //: /sn:0 {0}(210,96)(210,200){1}
//: {2}(208,202)(181,202)(181,220){3}
//: {4}(210,204)(210,221){5}
input G1;    //: /sn:0 {0}(512,91)(512,206){1}
//: {2}(514,208)(530,208)(530,220){3}
//: {4}(512,210)(512,219){5}
output O;    //: /sn:0 {0}(104,252)(104,281){1}
input Cin;    //: /sn:0 {0}(749,285)(737,285){1}
//: {2}(733,285)(712,285)(712,303){3}
//: {4}(735,287)(735,385)(721,385){5}
input G3;    //: /sn:0 {0}(186,96)(186,207){1}
//: {2}(188,209)(205,209)(205,221){3}
//: {4}(186,211)(186,220){5}
input P0;    //: /sn:0 {0}(685,89)(685,196){1}
//: {2}(683,198)(654,198)(654,217){3}
//: {4}(685,200)(685,217){5}
output S3;    //: /sn:0 /dp:1 {0}(248,308)(248,441){1}
input P2;    //: /sn:0 {0}(342,91)(342,197){1}
//: {2}(340,199)(315,199)(315,216){3}
//: {4}(342,201)(342,218){5}
output S2;    //: /sn:0 {0}(370,443)(370,307){1}
wire g1;    //: /sn:0 {0}(509,240)(509,360){1}
wire c0;    //: /sn:0 {0}(633,407)(633,417)(617,417)(617,283)(580,283)(580,291){1}
wire w51;    //: /sn:0 {0}(317,237)(317,360){1}
wire c1;    //: /sn:0 {0}(486,407)(486,416)(467,416)(467,275)(373,275)(373,286){1}
wire p3;    //: /sn:0 {0}(207,360)(207,280){1}
//: {2}(209,278)(246,278)(246,287){3}
//: {4}(207,276)(207,242){5}
wire p2;    //: /sn:0 {0}(339,360)(339,277){1}
//: {2}(341,275)(368,275)(368,286){3}
//: {4}(339,273)(339,239){5}
wire p1;    //: /sn:0 {0}(532,360)(532,285){1}
//: {2}(534,283)(575,283)(575,291){3}
//: {4}(532,281)(532,241){5}
wire w49;    //: /sn:0 {0}(656,238)(656,360){1}
wire p0;    //: /sn:0 {0}(682,360)(682,287){1}
//: {2}(684,285)(707,285)(707,303){3}
//: {4}(682,283)(682,238){5}
wire w2;    //: /sn:0 {0}(106,302)(106,322)(279,322){1}
//: {2}(281,320)(281,277)(251,277)(251,287){3}
//: {4}(281,324)(281,419)(302,419)(302,407){5}
wire w55;    //: /sn:0 {0}(183,241)(183,360){1}
//: enddecls

  //: input g8 (P2) @(342,89) /sn:0 /R:3 /w:[ 0 ]
  //: output g4 (S2) @(370,440) /sn:0 /R:3 /w:[ 0 ]
  //: joint g61 (P2) @(342, 199) /w:[ -1 1 2 4 ]
  //: input g13 (G3) @(186,94) /sn:0 /R:3 /w:[ 0 ]
  //: output g3 (S1) @(577,444) /sn:0 /R:3 /w:[ 0 ]
  CLA g55 (.G3(w55), .P3(p3), .G2(w51), .P2(p2), .G1(g1), .P1(p1), .G0(w49), .P0(p0), .Cin(Cin), .C3(C3), .Ps(Ps), .Gs(Gs), .C2(w2), .C1(c1), .C0(c0));   //: @(127, 361) /sz:(593, 45) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>1 Ti3>0 Ti4>1 Ti5>0 Ti6>1 Ti7>0 Ri0>5 Lo0<3 Bo0<1 Bo1<1 Bo2<5 Bo3<0 Bo4<0 ]
  //: output g2 (S0) @(696,444) /sn:0 /R:3 /w:[ 1 ]
  and g65 (.I0(G2), .I1(P2), .Z(w51));   //: @(317,227) /sn:0 /R:3 /w:[ 5 3 0 ]
  xor g76 (.I0(c0), .I1(p1), .Z(S1));   //: @(577,302) /sn:0 /R:3 /w:[ 1 3 1 ]
  xor g77 (.I0(c1), .I1(p2), .Z(S2));   //: @(370,297) /sn:0 /R:3 /w:[ 1 3 1 ]
  //: joint g59 (P3) @(210, 202) /w:[ -1 1 2 4 ]
  //: output g1 (Ps) @(206,438) /sn:0 /R:3 /w:[ 0 ]
  and g72 (.I0(G3), .I1(P3), .Z(w55));   //: @(183,231) /sn:0 /R:3 /w:[ 5 3 0 ]
  //: joint g64 (P0) @(685, 198) /w:[ -1 1 2 4 ]
  //: joint g16 (Cin) @(735, 285) /w:[ 1 -1 2 4 ]
  //: input g11 (G1) @(512,89) /sn:0 /R:3 /w:[ 0 ]
  //: input g10 (G0) @(659,88) /sn:0 /R:3 /w:[ 0 ]
  xor g78 (.I0(w2), .I1(p3), .Z(S3));   //: @(248,298) /sn:0 /R:3 /w:[ 3 3 0 ]
  //: joint g19 (C3) @(101, 381) /w:[ 2 4 1 -1 ]
  //: input g6 (P0) @(685,87) /sn:0 /R:3 /w:[ 0 ]
  xor g69 (.I0(P3), .I1(G3), .Z(p3));   //: @(207,232) /sn:0 /R:3 /w:[ 5 3 5 ]
  //: input g9 (P3) @(210,94) /sn:0 /R:3 /w:[ 0 ]
  //: input g7 (P1) @(535,88) /sn:0 /R:3 /w:[ 0 ]
  xor g57 (.I0(P0), .I1(G0), .Z(p0));   //: @(682,228) /sn:0 /R:3 /w:[ 5 3 5 ]
  //: joint g75 (G2) @(320, 204) /w:[ 2 1 -1 4 ]
  //: input g15 (Cin) @(751,285) /sn:0 /R:2 /w:[ 0 ]
  //: joint g71 (G1) @(512, 208) /w:[ 2 1 -1 4 ]
  //: output g20 (O) @(104,255) /sn:0 /R:1 /w:[ 0 ]
  //: joint g68 (P1) @(535, 201) /w:[ -1 1 2 4 ]
  and g62 (.I0(G0), .I1(P0), .Z(w49));   //: @(656,228) /sn:0 /R:3 /w:[ 5 3 0 ]
  //: joint g17 (w2) @(281, 322) /w:[ -1 2 1 4 ]
  and g63 (.I0(G1), .I1(P1), .Z(g1));   //: @(509,230) /sn:0 /R:3 /w:[ 5 3 0 ]
  //: joint g83 (p2) @(339, 275) /w:[ 2 4 -1 1 ]
  //: joint g74 (G0) @(659, 205) /w:[ 2 1 -1 4 ]
  //: output g14 (C3) @(82,381) /sn:0 /R:2 /w:[ 0 ]
  //: output g5 (S3) @(248,438) /sn:0 /R:3 /w:[ 1 ]
  xor g79 (.I0(Cin), .I1(p0), .Z(S0));   //: @(709,314) /sn:0 /R:3 /w:[ 3 3 0 ]
  //: joint g84 (p3) @(207, 278) /w:[ 2 4 -1 1 ]
  xor g60 (.I0(P1), .I1(G1), .Z(p1));   //: @(532,231) /sn:0 /R:3 /w:[ 5 3 5 ]
  //: joint g81 (p0) @(682, 285) /w:[ 2 4 -1 1 ]
  //: output g0 (Gs) @(188,439) /sn:0 /R:3 /w:[ 0 ]
  xor g70 (.I0(P2), .I1(G2), .Z(p2));   //: @(339,229) /sn:0 /R:3 /w:[ 5 3 5 ]
  //: joint g66 (G3) @(186, 209) /w:[ 2 1 -1 4 ]
  //: joint g82 (p1) @(532, 283) /w:[ 2 4 -1 1 ]
  //: input g12 (G2) @(320,89) /sn:0 /R:3 /w:[ 0 ]
  xor g18 (.I0(C3), .I1(w2), .Z(O));   //: @(104,291) /sn:0 /R:1 /w:[ 5 0 1 ]

endmodule

module ULA(ctrlULA, B, R, A, S);
//: interface  /sz:(40, 40) /bd:[ ]
supply0 w6;    //: /sn:0 /dp:1 {0}(571,688)(473,688){1}
//: {2}(471,686)(471,641){3}
//: {4}(473,639)(537,639){5}
//: {6}(471,637)(471,588){7}
//: {8}(473,586)(507,586){9}
//: {10}(471,584)(471,539)(483,539){11}
//: {12}(471,690)(471,735){13}
input [15:0] B;    //: /sn:0 /dp:1 {0}(52,501)(108,501)(108,264){1}
//: {2}(110,262)(255,262){3}
//: {4}(108,260)(108,201){5}
//: {6}(110,199)(255,199){7}
//: {8}(108,197)(108,122){9}
//: {10}(110,120)(255,120){11}
//: {12}(108,118)(108,49)(255,49){13}
input [15:0] A;    //: /sn:0 {0}(255,375)(81,375){1}
//: {2}(79,373)(79,314){3}
//: {4}(81,312)(255,312){5}
//: {6}(79,310)(79,234){7}
//: {8}(81,232)(255,232){9}
//: {10}(79,230)(79,164){11}
//: {12}(81,162)(255,162){13}
//: {14}(79,160)(79,90){15}
//: {16}(81,88)(255,88){17}
//: {18}(79,86)(79,17)(255,17){19}
//: {20}(79,377)(79,473)(52,473){21}
supply0 [15:0] w37;    //: /sn:0 {0}(637,349)(637,253){1}
//: {2}(639,251)(650,251){3}
//: {4}(637,249)(637,244)(650,244){5}
output [15:0] R;    //: /sn:0 /dp:1 {0}(679,255)(802,255){1}
supply0 [3:0] w11;    //: /sn:0 {0}(650,467)(611,467){1}
//: {2}(609,465)(609,460)(650,460){3}
//: {4}(607,467)(604,467)(604,494){5}
output [3:0] S;    //: /sn:0 {0}(806,471)(679,471){1}
input [2:0] ctrlULA;    //: /sn:0 /dp:3 {0}(711,-38)(711,414){1}
//: {2}(709,416)(666,416)(666,278){3}
//: {4}(711,418)(711,537)(666,537)(666,494){5}
wire z14;    //: /sn:0 /dp:1 {0}(507,566)(495,566)(495,264)(329,264){1}
wire w7;    //: /sn:0 /dp:1 {0}(329,127)(437,127)(437,460)(454,460){1}
wire w16;    //: /sn:0 /dp:1 {0}(329,99)(449,99)(449,490)(454,490){1}
wire z15;    //: /sn:0 /dp:1 {0}(537,619)(523,619)(523,330)(329,330){1}
wire w14;    //: /sn:0 /dp:1 {0}(507,576)(491,576)(491,273)(329,273){1}
wire w15;    //: /sn:0 /dp:1 {0}(329,108)(443,108)(443,480)(454,480){1}
wire z12;    //: /sn:0 {0}(329,192)(472,192)(472,519)(483,519){1}
wire p10;    //: /sn:0 /dp:1 {0}(574,445)(553,445)(553,47)(329,47){1}
wire [3:0] w19;    //: /sn:0 {0}(650,487)(632,487)(632,624)(543,624){1}
wire w3;    //: /sn:0 {0}(255,134)(194,134)(194,65){1}
//: {2}(196,63)(255,63){3}
//: {4}(194,61)(194,-37)(186,-37){5}
wire [3:0] w0;    //: /sn:0 {0}(650,447)(589,447)(589,440)(580,440){1}
wire n15;    //: /sn:0 {0}(329,322)(529,322)(529,609)(537,609){1}
wire [15:0] ressul;    //: /sn:0 {0}(329,16)(645,16)(645,231)(650,231){1}
wire p16;    //: /sn:0 /dp:1 {0}(571,678)(342,678)(342,416)(330,416){1}
wire z16;    //: /sn:0 /dp:1 {0}(571,668)(348,668)(348,408)(330,408){1}
wire n16;    //: /sn:0 {0}(330,400)(351,400)(351,658)(571,658){1}
wire [3:0] w20;    //: /sn:0 {0}(650,494)(640,494)(640,673)(577,673){1}
wire [15:0] w1;    //: /sn:0 {0}(650,264)(540,264)(540,232)(329,232){1}
wire p15;    //: /sn:0 /dp:1 {0}(537,629)(518,629)(518,339)(329,339){1}
wire n14;    //: /sn:0 {0}(329,252)(500,252)(500,556)(507,556){1}
wire z10;    //: /sn:0 /dp:1 {0}(574,435)(558,435)(558,37)(329,37){1}
wire w8;    //: /sn:0 /dp:1 {0}(329,118)(439,118)(439,470)(454,470){1}
wire [3:0] w18;    //: /sn:0 {0}(650,480)(624,480)(624,571)(513,571){1}
wire n10;    //: /sn:0 /dp:1 {0}(574,425)(563,425)(563,28)(329,28){1}
wire p13;    //: /sn:0 /dp:1 {0}(483,529)(468,529)(468,201)(329,201){1}
wire o10;    //: /sn:0 /dp:1 {0}(574,455)(548,455)(548,56)(329,56){1}
wire [15:0] w12;    //: /sn:0 /dp:1 {0}(650,271)(541,271)(541,304)(329,304){1}
wire [3:0] w10;    //: /sn:0 {0}(650,474)(622,474)(622,524)(489,524){1}
wire [15:0] R0;    //: /sn:0 {0}(330,373)(589,373)(589,278)(650,278){1}
wire n12;    //: /sn:0 /dp:1 {0}(483,509)(476,509)(476,182)(329,182){1}
wire [15:0] w13;    //: /sn:0 {0}(329,163)(588,163)(588,258)(650,258){1}
wire [3:0] w5;    //: /sn:0 /dp:1 {0}(650,454)(594,454)(594,475)(460,475){1}
wire [15:0] ressul0;    //: /sn:0 {0}(329,87)(636,87)(636,238)(650,238){1}
//: enddecls

  //: joint g4 (A) @(79, 88) /w:[ 16 18 -1 15 ]
  NOT g8 (.A(A), .p(p15), .z(z15), .n(n15), .R(w12));   //: @(256, 293) /sz:(72, 66) /sn:0 /p:[ Li0>5 Ro0<1 Ro1<1 Ro2<0 Ro3<1 ]
  //: joint g3 (w6) @(471, 586) /w:[ 8 10 -1 7 ]
  IDENTIDADE g37 (.A(A), .p(p16), .n(n16), .z(z16), .R(R0));   //: @(256, 361) /sz:(73, 66) /sn:0 /p:[ Li0>0 Ro0<1 Ro1<0 Ro2<1 Ro3<0 ]
  concat g13 (.I0(o10), .I1(p10), .I2(z10), .I3(n10), .Z(w0));   //: @(579,440) /sn:0 /w:[ 0 0 0 0 1 ] /dr:0
  //: input g2 (ctrlULA) @(711,-40) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (B) @(50,501) /sn:0 /w:[ 0 ]
  //: joint g11 (A) @(79, 375) /w:[ 1 2 -1 20 ]
  //: joint g16 (w37) @(637, 251) /w:[ 2 4 -1 1 ]
  concat g28 (.I0(w6), .I1(p15), .I2(z15), .I3(n15), .Z(w19));   //: @(542,624) /sn:0 /w:[ 5 0 0 1 1 ] /dr:0
  //: joint g10 (B) @(108, 262) /w:[ 2 4 -1 1 ]
  //: joint g27 (w6) @(471, 639) /w:[ 4 6 -1 3 ]
  //: joint g32 (A) @(79, 312) /w:[ 4 6 -1 3 ]
  //: joint g19 (ctrlULA) @(711, 416) /w:[ -1 1 2 4 ]
  AND g6 (.B(B), .A(A), .p(w14), .z(z14), .n(n14), .R(w1));   //: @(256, 216) /sz:(72, 75) /sn:0 /p:[ Li0>3 Li1>9 Ro0<1 Ro1<1 Ro2<0 Ro3<1 ]
  //: joint g9 (A) @(79, 232) /w:[ 8 10 -1 7 ]
  OR g7 (.B(B), .A(A), .z(z12), .p(p13), .n(n12), .R(w13));   //: @(256, 146) /sz:(72, 68) /sn:0 /p:[ Li0>7 Li1>13 Ro0<0 Ro1<1 Ro2<1 Ro3<0 ]
  //: joint g31 (A) @(79, 162) /w:[ 12 14 -1 11 ]
  concat g20 (.I0(w16), .I1(w15), .I2(w8), .I3(w7), .Z(w5));   //: @(459,475) /sn:0 /w:[ 1 1 1 1 1 ] /dr:0
  //: supply0 g15 (w37) @(637,355) /sn:0 /w:[ 0 ]
  ADD g29 (.Cin(w3), .B(B), .A(A), .o(o10), .p(p10), .z(z10), .n(n10), .R(ressul));   //: @(256, 5) /sz:(72, 68) /sn:0 /p:[ Li0>3 Li1>13 Li2>19 Ro0<1 Ro1<1 Ro2<1 Ro3<1 Ro4<0 ]
  concat g25 (.I0(w6), .I1(w14), .I2(z14), .I3(n14), .Z(w18));   //: @(512,571) /sn:0 /w:[ 9 0 0 1 1 ] /dr:0
  mux g17 (.I0(w0), .I1(w5), .I2(w11), .I3(w11), .I4(w10), .I5(w18), .I6(w19), .I7(w20), .S(ctrlULA), .Z(S));   //: @(666,471) /sn:0 /R:1 /w:[ 0 0 3 0 0 0 0 0 5 1 ] /ss:0 /do:0
  //: joint g5 (B) @(108, 120) /w:[ 10 12 -1 9 ]
  mux g14 (.I0(ressul), .I1(ressul0), .I2(w37), .I3(w37), .I4(w13), .I5(w1), .I6(w12), .I7(R0), .S(ctrlULA), .Z(R));   //: @(666,255) /sn:0 /R:1 /w:[ 1 1 5 3 1 0 0 1 3 0 ] /ss:0 /do:0
  //: joint g44 (B) @(108, 199) /w:[ 6 8 -1 5 ]
  concat g24 (.I0(w6), .I1(p13), .I2(z12), .I3(n12), .Z(w10));   //: @(488,524) /sn:0 /w:[ 11 0 1 0 1 ] /dr:0
  concat g36 (.I0(w6), .I1(p16), .I2(z16), .I3(n16), .Z(w20));   //: @(576,673) /sn:0 /w:[ 0 0 0 1 1 ] /dr:0
  //: supply0 g21 (w11) @(604,500) /sn:0 /w:[ 5 ]
  //: switch Cin (w3) @(169,-37) /w:[ 5 ] /st:0
  //: output g23 (R) @(799,255) /sn:0 /w:[ 1 ]
  //: joint g22 (w6) @(471, 688) /w:[ 1 2 -1 12 ]
  //: supply0 g26 (w6) @(471,741) /sn:0 /w:[ 13 ]
  //: input g0 (A) @(50,473) /sn:0 /w:[ 21 ]
  //: output g18 (S) @(803,471) /sn:0 /w:[ 0 ]
  //: joint g12 (w11) @(609, 467) /w:[ 1 2 4 -1 ]
  //: joint g33 (w3) @(194, 63) /w:[ 2 4 -1 1 ]
  SUB g30 (.Cin(w3), .B(B), .A(A), .o(w7), .p(w8), .z(w15), .n(w16), .R(ressul0));   //: @(256, 76) /sz:(72, 68) /sn:0 /p:[ Li0>0 Li1>11 Li2>17 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 ]

endmodule

module D4bitCLAAdder();
//: interface  /sz:(40, 40) /bd:[ ]
//: enddecls


endmodule

module SOMADOR();
//: interface  /sz:(40, 40) /bd:[ ]
//: enddecls


endmodule

module IDENTIDADE(n, p, R, A, z);
//: interface  /sz:(40, 40) /bd:[ ]
output p;    //: /sn:0 /dp:1 {0}(530,175)(555,175){1}
output z;    //: /sn:0 /dp:1 {0}(464,217)(497,217){1}
//: {2}(501,217)(555,217){3}
//: {4}(499,215)(499,177)(509,177){5}
input [15:0] A;    //: /sn:0 {0}(73,160)(141,160){1}
output [15:0] R;    //: /sn:0 /dp:1 {0}(517,83)(305,83)(305,158){1}
//: {2}(303,160)(230,160){3}
//: {4}(305,162)(305,219)(356,219){5}
output n;    //: /sn:0 /dp:3 {0}(362,144)(433,144){1}
//: {2}(435,142)(435,137)(498,137){3}
//: {4}(502,137)(554,137){5}
//: {6}(500,139)(500,172)(509,172){7}
//: {8}(435,146)(435,180)(443,180){9}
wire w7;    //: /sn:0 {0}(147,135)(224,135){1}
wire w56;    //: /sn:0 {0}(224,215)(147,215){1}
wire w14;    //: /sn:0 {0}(147,185)(224,185){1}
wire w16;    //: /sn:0 {0}(147,165)(224,165){1}
wire w19;    //: /sn:0 {0}(443,245)(427,245)(427,274)(362,274){1}
wire w4;    //: /sn:0 {0}(362,294)(435,294)(435,255)(443,255){1}
wire w15;    //: /sn:0 {0}(147,175)(224,175){1}
wire w3;    //: /sn:0 {0}(147,85)(224,85){1}
wire w34;    //: /sn:0 {0}(147,95)(224,95){1}
wire w21;    //: /sn:0 {0}(362,254)(416,254)(416,235)(443,235){1}
wire w31;    //: /sn:0 {0}(362,154)(432,154)(432,185)(443,185){1}
wire w28;    //: /sn:0 {0}(362,184)(422,184)(422,200)(443,200){1}
wire w24;    //: /sn:0 {0}(362,224)(402,224)(402,220)(443,220){1}
wire w23;    //: /sn:0 {0}(362,234)(408,234)(408,225)(443,225){1}
wire w20;    //: /sn:0 {0}(362,264)(421,264)(421,240)(443,240){1}
wire w1;    //: /sn:0 {0}(147,235)(183,235)(224,235){1}
wire w25;    //: /sn:0 {0}(147,145)(224,145){1}
wire w18;    //: /sn:0 {0}(362,284)(432,284)(432,250)(443,250){1}
wire w8;    //: /sn:0 {0}(147,125)(224,125){1}
wire w30;    //: /sn:0 {0}(362,164)(429,164)(429,190)(443,190){1}
wire w22;    //: /sn:0 {0}(362,244)(412,244)(412,230)(443,230){1}
wire w17;    //: /sn:0 {0}(147,155)(224,155){1}
wire w12;    //: /sn:0 {0}(147,205)(224,205){1}
wire w10;    //: /sn:0 {0}(147,115)(224,115){1}
wire w27;    //: /sn:0 {0}(362,194)(419,194)(419,205)(443,205){1}
wire w13;    //: /sn:0 {0}(147,195)(224,195){1}
wire w5;    //: /sn:0 {0}(147,225)(224,225){1}
wire w33;    //: /sn:0 {0}(147,105)(224,105){1}
wire w29;    //: /sn:0 {0}(362,174)(425,174)(425,195)(443,195){1}
wire w9;    //: /sn:0 {0}(443,215)(402,215)(402,214)(362,214){1}
wire w26;    //: /sn:0 {0}(362,204)(415,204)(415,210)(443,210){1}
//: enddecls

  //: joint g4 (z) @(499, 217) /w:[ 2 4 1 -1 ]
  //: output g8 (n) @(551,137) /sn:0 /w:[ 5 ]
  //: output g13 (p) @(552,175) /sn:0 /w:[ 1 ]
  //: output g3 (R) @(514,83) /sn:0 /w:[ 0 ]
  nor g2 (.I0(n), .I1(z), .Z(p));   //: @(520,175) /sn:0 /w:[ 7 5 0 ]
  //: joint g1 (n) @(435, 144) /w:[ -1 2 1 8 ]
  concat g11 (.I0(w4), .I1(w18), .I2(w19), .I3(w20), .I4(w21), .I5(w22), .I6(w23), .I7(w24), .I8(w9), .I9(w26), .I10(w27), .I11(w28), .I12(w29), .I13(w30), .I14(w31), .I15(n), .Z(R));   //: @(357,219) /sn:0 /R:2 /w:[ 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 5 ] /dr:1
  //: joint g6 (n) @(500, 137) /w:[ 4 -1 3 6 ]
  //: joint g7 (R) @(305, 160) /w:[ -1 1 2 4 ]
  concat g15 (.I0(w1), .I1(w5), .I2(w56), .I3(w12), .I4(w13), .I5(w14), .I6(w15), .I7(w16), .I8(w17), .I9(w25), .I10(w7), .I11(w8), .I12(w10), .I13(w33), .I14(w34), .I15(w3), .Z(A));   //: @(142,160) /sn:0 /R:2 /w:[ 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:1
  concat g17 (.I0(w1), .I1(w5), .I2(w56), .I3(w12), .I4(w13), .I5(w14), .I6(w15), .I7(w16), .I8(w17), .I9(w25), .I10(w7), .I11(w8), .I12(w10), .I13(w33), .I14(w34), .I15(w3), .Z(R));   //: @(229,160) /sn:0 /w:[ 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 3 ] /dr:0
  nor g5 (.I0(n), .I1(w31), .I2(w30), .I3(w29), .I4(w28), .I5(w27), .I6(w26), .I7(w9), .I8(w24), .I9(w23), .I10(w22), .I11(w21), .I12(w20), .I13(w19), .I14(w18), .I15(w4), .Z(z));   //: @(454,217) /sn:0 /w:[ 9 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 ]
  //: input g0 (A) @(71,160) /sn:0 /w:[ 0 ]
  //: output g12 (z) @(552,217) /sn:0 /w:[ 3 ]

endmodule

module main;    //: root_module
wire p;    //: /sn:0 {0}(657,322)(657,351){1}
wire [15:0] B;    //: /sn:0 /dp:1 {0}(461,246)(505,246){1}
wire z;    //: /sn:0 {0}(642,322)(642,351){1}
wire LoadReg;    //: /sn:0 {0}(204,108)(291,108)(291,131){1}
wire [15:0] A;    //: /sn:0 /dp:1 {0}(368,199)(505,199){1}
wire w0;    //: /sn:0 {0}(437,424)(448,424)(448,269){1}
wire [4:0] w3;    //: /sn:0 /dp:1 {0}(185,402)(185,419)(265,419){1}
wire [3:0] RBA;    //: /sn:0 /dp:1 {0}(185,290)(185,301)(237,301)(237,324)(264,324){1}
wire en;    //: /sn:0 /dp:1 {0}(601,307)(589,307)(589,419)(581,419){1}
wire [15:0] R;    //: /sn:0 /dp:3 {0}(589,83)(589,105){1}
//: {2}(587,107)(327,107)(327,131){3}
//: {4}(589,109)(589,233){5}
//: {6}(591,235)(659,235)(659,181){7}
//: {8}(587,235)(570,235){9}
wire [15:0] DataOutBusB;    //: /sn:0 /dp:1 {0}(368,236)(432,236){1}
wire o;    //: /sn:0 {0}(672,322)(672,351){1}
wire [15:0] Imm;    //: /sn:0 /dp:1 {0}(367,418)(386,418)(386,256)(432,256){1}
wire CLK;    //: /sn:0 /dp:1 {0}(712,303)(726,303)(726,463)(237,463){1}
//: {2}(235,461)(235,387)(264,387){3}
//: {4}(233,463)(147,463){5}
wire [3:0] RD;    //: /sn:0 /dp:1 {0}(186,231)(186,244)(238,244)(238,277)(264,277){1}
wire Reset;    //: /sn:0 /dp:1 {0}(264,171)(203,171){1}
wire n;    //: /sn:0 {0}(627,322)(627,351){1}
wire [3:0] RBB;    //: /sn:0 {0}(264,355)(186,355)(186,338){1}
wire [2:0] w5;    //: /sn:0 {0}(494,409)(494,320)(505,320){1}
wire [3:0] S;    //: /sn:0 /dp:1 {0}(601,289)(570,289){1}
//: enddecls

  led g4 (.I(z));   //: @(642,358) /sn:0 /R:2 /w:[ 1 ] /type:0
  REGSTAT g8 (.en(en), .S(S), .CLK(CLK), .o(o), .p(p), .z(z), .n(n));   //: @(602, 280) /sz:(109, 41) /sn:0 /p:[ Li0>0 Li1>0 Ri0>0 Bo0<0 Bo1<0 Bo2<0 Bo3<0 ]
  Extensao_Sinal g3 (.Imm5(w3), .Imm16(Imm));   //: @(266, 412) /sz:(100, 41) /sn:0 /p:[ Li0>1 Ro0<0 ]
  //: joint g13 (CLK) @(235, 463) /w:[ 1 2 4 -1 ]
  REGISTRADORES g2 (.LoadReg(LoadReg), .R(R), .Reset(Reset), .CLK(CLK), .RegDst(RD), .RegBusB(RBB), .RegBusA(RBA), .DataOutBusA(A), .DataOutBusB(DataOutBusB));   //: @(265, 132) /sz:(102, 268) /sn:0 /p:[ Ti0>1 Ti1>3 Li0>0 Li1>3 Li2>1 Li3>0 Li4>1 Ro0<0 Ro1<0 ]
  mux g1 (.I0(Imm), .I1(DataOutBusB), .S(w0), .Z(B));   //: @(448,246) /sn:0 /R:1 /w:[ 1 1 1 0 ] /ss:0 /do:0
  //: dip RegB (RBB) @(186,328) /w:[ 1 ] /st:0
  //: switch LoadReg (LoadReg) @(187,108) /w:[ 0 ] /st:1
  led g11 (.I(R));   //: @(659,174) /sn:0 /w:[ 7 ] /type:3
  clock g10 (.Z(CLK));   //: @(134,463) /sn:0 /w:[ 5 ] /omega:500 /phi:0 /duty:80
  led g6 (.I(p));   //: @(657,358) /sn:0 /R:2 /w:[ 1 ] /type:0
  led g7 (.I(n));   //: @(627,358) /sn:0 /R:2 /w:[ 1 ] /type:0
  led g9 (.I(o));   //: @(672,358) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: dip Imm5 (w3) @(185,392) /w:[ 0 ] /st:31
  //: dip RegA (RBA) @(185,280) /w:[ 0 ] /st:0
  ULA ULA (.ctrlULA(w5), .B(B), .A(A), .R(R), .S(S));   //: @(506, 147) /sz:(63, 191) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Ro0<9 Ro1<1 ]
  //: switch En (en) @(564,419) /w:[ 1 ] /st:0
  //: dip RegDst (RD) @(186,221) /w:[ 0 ] /st:0
  led g5 (.I(R));   //: @(589,76) /sn:0 /w:[ 0 ] /type:1
  //: switch Reset (Reset) @(186,171) /w:[ 1 ] /st:0
  //: joint g0 (R) @(589, 235) /w:[ 6 5 8 -1 ]
  //: joint g12 (R) @(589, 107) /w:[ -1 1 2 4 ]
  //: switch SelB (w0) @(420,424) /w:[ 0 ] /st:0
  //: dip ctrlULA (w5) @(494,420) /R:2 /w:[ 0 ] /st:0

endmodule

module Extensao_Sinal(Imm16, Imm5);
//: interface  /sz:(40, 40) /bd:[ ]
input [4:0] Imm5;    //: /sn:0 {0}(214,214)(130,214){1}
output [15:0] Imm16;    //: /sn:0 /dp:1 {0}(436,322)(436,345)(479,345){1}
wire w7;    //: /sn:0 {0}(401,316)(401,250){1}
//: {2}(403,248)(419,248){3}
//: {4}(423,248)(439,248){5}
//: {6}(443,248)(459,248){7}
//: {8}(463,248)(479,248){9}
//: {10}(483,248)(501,248)(501,316){11}
//: {12}(481,250)(481,316){13}
//: {14}(461,250)(461,316){15}
//: {16}(441,250)(441,316){17}
//: {18}(421,250)(421,316){19}
//: {20}(401,246)(401,236){21}
//: {22}(403,234)(409,234){23}
//: {24}(413,234)(429,234){25}
//: {26}(433,234)(449,234){27}
//: {28}(453,234)(469,234){29}
//: {30}(473,234)(489,234){31}
//: {32}(493,234)(511,234)(511,316){33}
//: {34}(491,236)(491,316){35}
//: {36}(471,236)(471,316){37}
//: {38}(451,236)(451,316){39}
//: {40}(431,236)(431,316){41}
//: {42}(411,236)(411,316){43}
//: {44}(399,234)(220,234){45}
wire w0;    //: /sn:0 /dp:1 {0}(371,316)(371,269)(326,269)(326,204)(220,204){1}
wire w3;    //: /sn:0 {0}(220,194)(313,194)(313,277)(361,277)(361,316){1}
wire w8;    //: /sn:0 {0}(220,214)(340,214)(340,260)(381,260)(381,316){1}
wire w9;    //: /sn:0 {0}(220,224)(353,224)(353,248)(391,248)(391,316){1}
//: enddecls

  //: joint g8 (w7) @(411, 234) /w:[ 24 -1 23 42 ]
  //: joint g4 (w7) @(491, 234) /w:[ 32 -1 31 34 ]
  //: joint g13 (w7) @(401, 248) /w:[ 2 20 -1 1 ]
  concat g3 (.I0(w3), .I1(w0), .I2(w8), .I3(w9), .I4(w7), .Z(Imm5));   //: @(215,214) /sn:0 /R:2 /w:[ 0 1 0 0 45 0 ] /dr:0
  concat g2 (.I0(w3), .I1(w0), .I2(w8), .I3(w9), .I4(w7), .I5(w7), .I6(w7), .I7(w7), .I8(w7), .I9(w7), .I10(w7), .I11(w7), .I12(w7), .I13(w7), .I14(w7), .I15(w7), .Z(Imm16));   //: @(436,321) /sn:0 /R:3 /w:[ 1 0 1 1 0 43 19 41 17 39 15 37 13 35 11 33 0 ] /dr:0
  //: output g1 (Imm16) @(476,345) /sn:0 /w:[ 1 ]
  //: joint g11 (w7) @(421, 248) /w:[ 4 -1 3 18 ]
  //: joint g10 (w7) @(441, 248) /w:[ 6 -1 5 16 ]
  //: joint g6 (w7) @(451, 234) /w:[ 28 -1 27 38 ]
  //: joint g9 (w7) @(461, 248) /w:[ 8 -1 7 14 ]
  //: joint g7 (w7) @(431, 234) /w:[ 26 -1 25 40 ]
  //: joint g14 (w7) @(481, 248) /w:[ 10 -1 9 12 ]
  //: joint g5 (w7) @(471, 234) /w:[ 30 -1 29 36 ]
  //: input g0 (Imm5) @(128,214) /sn:0 /w:[ 1 ]
  //: joint g12 (w7) @(401, 234) /w:[ 22 -1 44 21 ]

endmodule

module NOT(n, p, R, A, z);
//: interface  /sz:(40, 40) /bd:[ ]
output p;    //: /sn:0 {0}(512,197)(558,197){1}
output z;    //: /sn:0 /dp:1 {0}(452,239)(484,239){1}
//: {2}(488,239)(558,239){3}
//: {4}(486,237)(486,199)(491,199){5}
input [15:0] A;    //: /sn:0 {0}(104,241)(163,241){1}
output [15:0] R;    //: /sn:0 {0}(179,241)(263,241){1}
//: {2}(267,241)(344,241){3}
//: {4}(265,239)(265,105)(505,105){5}
output n;    //: /sn:0 /dp:3 {0}(350,166)(421,166){1}
//: {2}(423,164)(423,159)(482,159){3}
//: {4}(486,159)(556,159){5}
//: {6}(484,161)(484,194)(491,194){7}
//: {8}(423,168)(423,202)(431,202){9}
wire w4;    //: /sn:0 {0}(350,316)(423,316)(423,277)(431,277){1}
wire w19;    //: /sn:0 {0}(431,267)(415,267)(415,296)(350,296){1}
wire w21;    //: /sn:0 {0}(350,276)(404,276)(404,257)(431,257){1}
wire w31;    //: /sn:0 {0}(350,176)(420,176)(420,207)(431,207){1}
wire w28;    //: /sn:0 {0}(350,206)(410,206)(410,222)(431,222){1}
wire w20;    //: /sn:0 {0}(350,286)(409,286)(409,262)(431,262){1}
wire w23;    //: /sn:0 {0}(350,256)(396,256)(396,247)(431,247){1}
wire w24;    //: /sn:0 {0}(350,246)(390,246)(390,242)(431,242){1}
wire w18;    //: /sn:0 {0}(350,306)(420,306)(420,272)(431,272){1}
wire w30;    //: /sn:0 {0}(350,186)(417,186)(417,212)(431,212){1}
wire w22;    //: /sn:0 {0}(350,266)(400,266)(400,252)(431,252){1}
wire w27;    //: /sn:0 {0}(350,216)(407,216)(407,227)(431,227){1}
wire w29;    //: /sn:0 {0}(350,196)(413,196)(413,217)(431,217){1}
wire w9;    //: /sn:0 {0}(431,237)(390,237)(390,236)(350,236){1}
wire w26;    //: /sn:0 {0}(350,226)(403,226)(403,232)(431,232){1}
//: enddecls

  nor g4 (.I0(n), .I1(z), .Z(p));   //: @(502,197) /sn:0 /w:[ 7 5 0 ]
  //: output g8 (n) @(553,159) /sn:0 /w:[ 5 ]
  //: output g13 (p) @(555,197) /sn:0 /w:[ 1 ]
  //: output g3 (R) @(502,105) /sn:0 /w:[ 5 ]
  //: joint g2 (R) @(265, 241) /w:[ 2 4 1 -1 ]
  //: joint g1 (n) @(423, 166) /w:[ -1 2 1 8 ]
  concat g11 (.I0(w4), .I1(w18), .I2(w19), .I3(w20), .I4(w21), .I5(w22), .I6(w23), .I7(w24), .I8(w9), .I9(w26), .I10(w27), .I11(w28), .I12(w29), .I13(w30), .I14(w31), .I15(n), .Z(R));   //: @(345,241) /sn:0 /R:2 /w:[ 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 3 ] /dr:1
  //: joint g6 (n) @(484, 159) /w:[ 4 -1 3 6 ]
  //: joint g9 (z) @(486, 239) /w:[ 2 4 1 -1 ]
  not g7 (.I(A), .Z(R));   //: @(169,241) /sn:0 /w:[ 1 0 ]
  nor g5 (.I0(n), .I1(w31), .I2(w30), .I3(w29), .I4(w28), .I5(w27), .I6(w26), .I7(w9), .I8(w24), .I9(w23), .I10(w22), .I11(w21), .I12(w20), .I13(w19), .I14(w18), .I15(w4), .Z(z));   //: @(442,239) /sn:0 /w:[ 9 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 ]
  //: input g0 (A) @(102,241) /sn:0 /w:[ 0 ]
  //: output g12 (z) @(555,239) /sn:0 /w:[ 3 ]

endmodule

module ADD(B, A, Cin, n, R, o, z, p);
//: interface  /sz:(40, 40) /bd:[ ]
output p;    //: /sn:0 {0}(520,380)(491,380){1}
output z;    //: /sn:0 {0}(519,402)(450,402){1}
//: {2}(448,400)(448,382)(470,382){3}
//: {4}(446,402)(419,402){5}
input [15:0] B;    //: /sn:0 {0}(21,-350)(21,-405){1}
input [15:0] A;    //: /sn:0 {0}(592,-372)(592,-397){1}
output [15:0] R;    //: /sn:0 {0}(398,402)(344,402){1}
//: {2}(342,400)(342,373){3}
//: {4}(342,404)(342,426){5}
output o;    //: /sn:0 {0}(522,451)(-489,451)(-489,6)(-405,6){1}
input Cin;    //: /sn:0 {0}(942,-8)(977,-8){1}
//: {2}(981,-8)(995,-8){3}
//: {4}(979,-6)(979,90)(955,90){5}
output n;    //: /sn:0 {0}(521,343)(450,343){1}
//: {2}(446,343)(419,343){3}
//: {4}(415,343)(-194,343)(-194,29){5}
//: {6}(417,345)(417,367){7}
//: {8}(448,345)(448,377)(470,377){9}
wire w32;    //: /sn:0 {0}(31,28)(31,64){1}
wire w6;    //: /sn:0 {0}(766,-31)(766,-318)(76,-318)(76,-344){1}
wire w7;    //: /sn:0 {0}(424,-30)(424,-87)(536,-87)(536,-276)(36,-276)(36,-344){1}
wire c6;    //: /sn:0 {0}(632,112)(632,140)(617,140)(617,-7)(600,-7){1}
wire Ps;    //: /sn:0 {0}(-229,112)(-229,144)(-251,144)(-251,133){1}
wire p6;    //: /sn:0 {0}(390,64)(390,28){1}
wire w16;    //: /sn:0 {0}(607,-366)(607,-83)(529,-83)(529,-65)(435,-65)(435,-30){1}
wire a2;    //: /sn:0 {0}(777,-31)(777,-347)(647,-347)(647,-366){1}
wire w4;    //: /sn:0 {0}(287,367)(287,176)(894,176)(894,27){1}
wire w15;    //: /sn:0 {0}(617,-366)(617,-71)(539,-71)(539,-35)(501,-35)(501,-30){1}
wire b2;    //: /sn:0 {0}(843,-31)(843,-351)(657,-351)(657,-366){1}
wire w38;    //: /sn:0 {0}(227,28)(227,249)(347,249)(347,367){1}
wire w51;    //: /sn:0 {0}(-4,-344)(-4,-41)(65,-41)(65,-30){1}
wire w69;    //: /sn:0 {0}(702,64)(702,27){1}
wire a7;    //: /sn:0 {0}(-180,-29)(-180,-223)(547,-223)(547,-366){1}
wire a4;    //: /sn:0 {0}(76,-30)(76,-66)(173,-66)(173,-210)(567,-210)(567,-366){1}
wire w3;    //: /sn:0 {0}(-447,56)(-447,86)(-411,86){1}
wire b11;    //: /sn:0 {0}(142,-30)(142,-45)(182,-45)(182,-201)(577,-201)(577,-366){1}
wire w0;    //: /sn:0 {0}(-454,-85)(-454,-11)(-405,-11){1}
wire w66;    //: /sn:0 {0}(-143,29)(-143,301)(387,301)(387,367){1}
wire w64;    //: /sn:0 {0}(-359,-29)(-359,-247)(517,-247)(517,-366){1}
wire w34;    //: /sn:0 {0}(176,28)(176,280)(377,280)(377,367){1}
wire w63;    //: /sn:0 {0}(11,-30)(11,-70)(163,-70)(163,-218)(557,-218)(557,-366){1}
wire w54;    //: /sn:0 {0}(-34,-344)(-34,-267)(-240,-267)(-240,-29){1}
wire b3;    //: /sn:0 {0}(831,-31)(831,-325)(86,-325)(86,-344){1}
wire w58;    //: /sn:0 {0}(-177,29)(-177,327)(407,327)(407,367){1}
wire w28;    //: /sn:0 {0}(327,367)(327,224)(552,224)(552,28){1}
wire b6;    //: /sn:0 {0}(489,-30)(489,-95)(551,-95)(551,-285)(46,-285)(46,-344){1}
wire w36;    //: /sn:0 {0}(210,28)(210,258)(357,258)(357,367){1}
wire w20;    //: /sn:0 {0}(928,27)(928,154)(267,154)(267,367){1}
wire w23;    //: /sn:0 {0}(587,-366)(587,-192)(190,-192)(190,-30){1}
wire w1;    //: /sn:0 {0}(298,-17)(298,-4)(324,-4){1}
wire Gs;    //: /sn:0 {0}(-270,112)(-270,145)(-292,145)(-292,134){1}
wire b15;    //: /sn:0 {0}(-228,-29)(-228,-231)(537,-231)(537,-366){1}
wire w65;    //: /sn:0 {0}(-160,29)(-160,313)(397,313)(397,367){1}
wire a6;    //: /sn:0 {0}(-294,-29)(-294,-241)(527,-241)(527,-366){1}
wire a1;    //: /sn:0 {0}(549,-30)(549,-61)(627,-61)(627,-366){1}
wire w35;    //: /sn:0 {0}(193,28)(193,268)(367,268)(367,367){1}
wire w40;    //: /sn:0 {0}(-369,29)(-369,64){1}
wire w8;    //: /sn:0 {0}(297,367)(297,188)(877,188)(877,27){1}
wire b1;    //: /sn:0 {0}(878,-31)(878,-331)(96,-331)(96,-344){1}
wire w30;    //: /sn:0 {0}(337,367)(337,236)(535,236)(535,28){1}
wire b4;    //: /sn:0 {0}(687,-31)(687,-311)(66,-311)(66,-344){1}
wire w22;    //: /sn:0 {0}(597,-366)(597,-94)(518,-94)(518,-66)(370,-66)(370,-30){1}
wire a0;    //: /sn:0 {0}(891,-31)(891,-356)(667,-356)(667,-366){1}
wire w59;    //: /sn:0 {0}(712,-31)(712,-342)(637,-342)(637,-366){1}
wire b16;    //: /sn:0 {0}(-193,-29)(-193,-261)(-24,-261)(-24,-344){1}
wire w49;    //: /sn:0 {0}(16,-344)(16,-59)(177,-59)(177,-30){1}
wire cin2;    //: /sn:0 {0}(-129,-6)(-110,-6)(-110,124)(-96,124)(-96,112){1}
wire w2;    //: /sn:0 {0}(277,367)(277,165)(911,165)(911,27){1}
wire w11;    //: /sn:0 {0}(-62,-34)(-62,-14)(-35,-14){1}
wire w12;    //: /sn:0 {0}(644,-22)(644,-5)(666,-5){1}
wire b8;    //: /sn:0 {0}(536,-30)(536,-103)(563,-103)(563,-296)(56,-296)(56,-344){1}
wire w10;    //: /sn:0 {0}(307,367)(307,201)(586,201)(586,28){1}
wire w13;    //: /sn:0 {0}(317,367)(317,213)(569,213)(569,28){1}
wire w52;    //: /sn:0 {0}(-14,-344)(-14,-30){1}
wire w5;    //: /sn:0 {0}(360,64)(360,28){1}
wire p7;    //: /sn:0 {0}(732,64)(732,27){1}
wire w29;    //: /sn:0 {0}(1,28)(1,64){1}
wire p4;    //: /sn:0 {0}(-339,64)(-339,29){1}
wire w50;    //: /sn:0 {0}(6,-344)(6,-47)(130,-47)(130,-30){1}
wire w9;    //: /sn:0 {0}(-305,-29)(-305,-254)(-44,-254)(-44,-344){1}
wire c5;    //: /sn:0 {0}(267,112)(267,122)(254,122)(254,-7)(241,-7){1}
wire b5;    //: /sn:0 {0}(345,-30)(345,-267)(26,-267)(26,-344){1}
wire b13;    //: /sn:0 {0}(-384,-29)(-384,-279)(-54,-279)(-54,-344){1}
//: enddecls

  concat g4 (.I0(a0), .I1(b2), .I2(a2), .I3(w59), .I4(a1), .I5(w15), .I6(w16), .I7(w22), .I8(w23), .I9(b11), .I10(a4), .I11(w63), .I12(a7), .I13(b15), .I14(a6), .I15(w64), .Z(A));   //: @(592,-371) /sn:0 /R:1 /w:[ 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 ] /dr:0
  led g8 (.I(w0));   //: @(-454,-92) /sn:0 /w:[ 0 ] /type:0
  //: input g3 (B) @(21,-407) /sn:0 /R:3 /w:[ 1 ]
  led g13 (.I(w12));   //: @(644,-29) /sn:0 /w:[ 0 ] /type:0
  //: input g2 (A) @(592,-399) /sn:0 /R:3 /w:[ 1 ]
  //: input g1 (Cin) @(997,-8) /sn:0 /R:2 /w:[ 3 ]
  //: output g16 (n) @(518,343) /sn:0 /w:[ 0 ]
  led g11 (.I(w11));   //: @(-62,-41) /sn:0 /w:[ 0 ] /type:0
  //: joint g28 (z) @(448, 402) /w:[ 1 2 4 -1 ]
  Somador_CLA_4Bits g10 (.G3(b4), .G2(w6), .G1(b3), .P2(a2), .P3(w59), .P1(b2), .G0(b1), .P0(a0), .Cin(Cin), .C3(w12), .Gs(w69), .Ps(p7), .S3(w8), .S2(w4), .S1(w2), .S0(w20));   //: @(667, -30) /sz:(274, 56) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Bo2<1 Bo3<1 Bo4<1 Bo5<0 ]
  //: joint g27 (n) @(448, 343) /w:[ 1 -1 2 8 ]
  Somador_CLA_4Bits g19 (.G3(b13), .G2(w9), .G1(w54), .P2(a6), .P3(w64), .P1(b15), .G0(b16), .P0(a7), .Cin(cin2), .O(o), .C3(w0), .Gs(w40), .Ps(p4), .S3(n), .S2(w58), .S1(w65), .S0(w66));   //: @(-404, -28) /sz:(274, 56) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Ti3>0 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>0 Lo0<1 Lo1<1 Bo0<0 Bo1<1 Bo2<5 Bo3<0 Bo4<0 Bo5<0 ]
  concat g6 (.I0(w20), .I1(w2), .I2(w4), .I3(w8), .I4(w10), .I5(w13), .I6(w28), .I7(w30), .I8(w38), .I9(w36), .I10(w35), .I11(w34), .I12(w66), .I13(w65), .I14(w58), .I15(n), .Z(R));   //: @(342,372) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 7 3 ] /dr:0
  //: output g7 (R) @(342,423) /sn:0 /R:3 /w:[ 5 ]
  led g9 (.I(w3));   //: @(-447,49) /sn:0 /w:[ 0 ] /type:0
  //: joint g20 (R) @(342, 402) /w:[ 1 2 -1 4 ]
  //: joint g15 (n) @(417, 343) /w:[ 3 -1 4 6 ]
  //: output g29 (o) @(519,451) /sn:0 /w:[ 0 ]
  nor g25 (.I0(n), .I1(z), .Z(p));   //: @(481,380) /sn:0 /w:[ 9 3 1 ]
  Somador_CLA_4Bits g17 (.G3(b5), .G2(w7), .G1(b6), .P2(w16), .P3(w22), .P1(w15), .G0(b8), .P0(a1), .Cin(c6), .C3(w1), .Gs(w5), .Ps(p6), .S3(w30), .S2(w28), .S1(w13), .S0(w10));   //: @(325, -29) /sz:(274, 56) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>1 Ti4>1 Ti5>1 Ti6>0 Ti7>0 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Bo2<1 Bo3<1 Bo4<1 Bo5<1 ]
  concat g5 (.I0(b1), .I1(b3), .I2(w6), .I3(b4), .I4(b8), .I5(b6), .I6(w7), .I7(b5), .I8(w49), .I9(w50), .I10(w51), .I11(w52), .I12(b16), .I13(w54), .I14(w9), .I15(b13), .Z(B));   //: @(21,-349) /sn:0 /R:1 /w:[ 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 ] /dr:0
  //: output g24 (z) @(516,402) /sn:0 /w:[ 0 ]
  led g21 (.I(Ps));   //: @(-251,126) /sn:0 /w:[ 1 ] /type:0
  nor g23 (.I0(R), .Z(z));   //: @(409,402) /sn:0 /w:[ 0 5 ]
  //: output g26 (p) @(517,380) /sn:0 /w:[ 0 ]
  //: joint g0 (Cin) @(979, -8) /w:[ 2 -1 1 4 ]
  led g22 (.I(Gs));   //: @(-292,127) /sn:0 /w:[ 1 ] /type:0
  Somador_CLA_4Bits g18 (.G3(w52), .G2(w51), .G1(w50), .P2(a4), .P3(w63), .P1(b11), .G0(w49), .P0(w23), .Cin(c5), .C3(w11), .Gs(w29), .Ps(w32), .S3(w34), .S2(w35), .S1(w36), .S0(w38));   //: @(-34, -29) /sz:(274, 56) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>0 Ti4>0 Ti5>0 Ti6>1 Ti7>1 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Bo2<0 Bo3<0 Bo4<0 Bo5<0 ]
  led g12 (.I(w1));   //: @(298,-24) /sn:0 /w:[ 0 ] /type:0
  CLA g91 (.G3(w40), .P3(p4), .G2(w29), .P2(w32), .G1(w5), .P1(p6), .G0(w69), .P0(p7), .Cin(Cin), .C3(w3), .Ps(Ps), .Gs(Gs), .C2(cin2), .C1(c5), .C0(c6));   //: @(-410, 65) /sz:(1364, 46) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>1 Ti3>1 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>5 Lo0<1 Bo0<0 Bo1<0 Bo2<1 Bo3<0 Bo4<0 ]

endmodule

module CLA(C3, G1, P2, Ps, G0, G3, P1, C2, P0, P3, C1, C0, Cin, Gs, G2);
//: interface  /sz:(40, 40) /bd:[ ]
input G2;    //: /sn:0 /dp:1 {0}(372,282)(372,276)(337,276)(337,116){1}
//: {2}(337,112)(337,94){3}
//: {4}(335,114)(200,114)(200,226){5}
output Ps;    //: /sn:0 {0}(279,369)(279,345){1}
//: {2}(279,341)(279,247){3}
//: {4}(277,343)(141,343){5}
output C0;    //: /sn:0 {0}(621,371)(621,306){1}
input P1;    //: /sn:0 /dp:15 {0}(402,225)(402,182){1}
//: {2}(404,180)(503,180){3}
//: {4}(505,178)(505,96){5}
//: {6}(505,182)(505,228){7}
//: {8}(400,180)(383,180){9}
//: {10}(379,180)(283,180){11}
//: {12}(279,180)(250,180)(250,226){13}
//: {14}(281,182)(281,226){15}
//: {16}(381,182)(381,225){17}
output C3;    //: /sn:0 {0}(48,325)(74,325){1}
input G0;    //: /sn:0 {0}(386,225)(386,196)(508,196){1}
//: {2}(512,196)(617,196){3}
//: {4}(619,194)(619,102)(618,102)(618,100){5}
//: {6}(619,198)(619,285){7}
//: {8}(510,198)(510,228){9}
output C2;    //: /sn:0 /dp:1 {0}(380,371)(380,303){1}
output Gs;    //: /sn:0 {0}(227,368)(227,325){1}
//: {2}(227,321)(227,302){3}
//: {4}(225,323)(95,323){5}
input P3;    //: /sn:0 {0}(271,226)(271,164)(242,164){1}
//: {2}(238,164)(217,164){3}
//: {4}(213,164)(197,164){5}
//: {6}(195,162)(195,95){7}
//: {8}(195,166)(195,226){9}
//: {10}(215,166)(215,226){11}
//: {12}(240,166)(240,226){13}
input G1;    //: /sn:0 /dp:1 {0}(531,230)(531,218)(489,218){1}
//: {2}(487,216)(487,177){3}
//: {4}(487,173)(487,96){5}
//: {6}(485,175)(364,175){7}
//: {8}(360,175)(257,175){9}
//: {10}(253,175)(225,175)(225,226){11}
//: {12}(255,177)(255,226){13}
//: {14}(362,177)(362,203)(361,203)(361,226){15}
//: {16}(487,220)(487,277)(515,277)(515,281){17}
input Cin;    //: /sn:0 {0}(732,203)(651,203){1}
//: {2}(647,203)(543,203){3}
//: {4}(539,203)(414,203){5}
//: {6}(410,203)(155,203)(155,338)(141,338){7}
//: {8}(412,205)(412,225){9}
//: {10}(541,205)(541,230){11}
//: {12}(649,205)(649,226){13}
input G3;    //: /sn:0 /dp:1 {0}(219,281)(219,273)(177,273)(177,94){1}
input P0;    //: /sn:0 {0}(644,101)(644,184){1}
//: {2}(642,186)(538,186){3}
//: {4}(534,186)(409,186){5}
//: {6}(407,184)(407,174){7}
//: {8}(405,186)(286,186)(286,226){9}
//: {10}(407,188)(407,225){11}
//: {12}(536,188)(536,230){13}
//: {14}(644,188)(644,226){15}
output C1;    //: /sn:0 /dp:1 {0}(520,372)(520,302){1}
input P2;    //: /sn:0 {0}(220,226)(220,187)(243,187){1}
//: {2}(247,187)(274,187){3}
//: {4}(278,187)(354,187){5}
//: {6}(358,187)(374,187){7}
//: {8}(378,187)(397,187)(397,225){9}
//: {10}(376,189)(376,225){11}
//: {12}(356,185)(356,94){13}
//: {14}(356,189)(356,226){15}
//: {16}(276,189)(276,226){17}
//: {18}(245,189)(245,226){19}
wire w14;    //: /sn:0 {0}(405,246)(405,272)(387,272)(387,282){1}
wire w37;    //: /sn:0 /dp:1 {0}(520,281)(520,266)(507,266)(507,249){1}
wire w21;    //: /sn:0 {0}(224,281)(224,263)(197,263)(197,247){1}
wire w23;    //: /sn:0 {0}(377,282)(377,251)(358,251)(358,247){1}
wire w36;    //: /sn:0 /dp:1 {0}(525,281)(525,266)(536,266)(536,251){1}
wire w8;    //: /sn:0 {0}(248,247)(248,260)(234,260)(234,281){1}
wire w17;    //: /sn:0 {0}(381,246)(381,272)(382,272)(382,282){1}
wire w11;    //: /sn:0 {0}(120,340)(105,340)(105,328)(95,328){1}
wire w5;    //: /sn:0 {0}(220,247)(220,258)(229,258)(229,281){1}
wire w29;    //: /sn:0 {0}(646,247)(646,275)(624,275)(624,285){1}
//: enddecls

  and g4 (.I0(Cin), .I1(P0), .I2(P1), .I3(P2), .Z(w14));   //: @(405,236) /sn:0 /R:3 /w:[ 9 11 0 9 0 ]
  and g8 (.I0(G0), .I1(P1), .Z(w37));   //: @(507,239) /sn:0 /R:3 /w:[ 9 7 1 ]
  //: joint g51 (G1) @(255, 175) /w:[ 9 -1 10 12 ]
  //: joint g55 (P1) @(281, 180) /w:[ 11 -1 12 14 ]
  //: joint g37 (Ps) @(279, 343) /w:[ -1 2 4 1 ]
  //: output g34 (C3) @(51,325) /sn:0 /R:2 /w:[ 0 ]
  and g3 (.I0(P0), .I1(P1), .I2(P2), .I3(P3), .Z(Ps));   //: @(279,237) /sn:0 /R:3 /w:[ 9 15 17 0 3 ]
  or g13 (.I0(w29), .I1(G0), .Z(C0));   //: @(621,296) /sn:0 /R:3 /w:[ 1 7 1 ]
  and g2 (.I0(G1), .I1(P1), .I2(P2), .I3(P3), .Z(w8));   //: @(248,237) /sn:0 /R:3 /w:[ 13 13 19 13 0 ]
  and g1 (.I0(G1), .I1(P2), .I2(P3), .Z(w5));   //: @(220,237) /sn:0 /R:3 /w:[ 11 0 11 0 ]
  or g11 (.I0(w14), .I1(w17), .I2(w23), .I3(G2), .Z(C2));   //: @(380,293) /sn:0 /R:3 /w:[ 1 1 0 0 1 ]
  //: input g16 (G1) @(487,94) /sn:0 /R:3 /w:[ 5 ]
  //: joint g50 (P0) @(407, 186) /w:[ 5 6 8 10 ]
  //: joint g28 (Cin) @(541, 203) /w:[ 3 -1 4 10 ]
  or g10 (.I0(w8), .I1(w5), .I2(w21), .I3(G3), .Z(Gs));   //: @(227,292) /sn:0 /R:3 /w:[ 1 1 0 0 3 ]
  and g32 (.I0(Ps), .I1(Cin), .Z(w11));   //: @(130,340) /sn:0 /R:2 /w:[ 5 7 0 ]
  //: joint g27 (Cin) @(649, 203) /w:[ 1 -1 2 12 ]
  //: input g19 (P2) @(356,92) /sn:0 /R:3 /w:[ 13 ]
  //: joint g38 (G2) @(337, 114) /w:[ -1 2 4 1 ]
  and g6 (.I0(G1), .I1(P2), .Z(w23));   //: @(358,237) /sn:0 /R:3 /w:[ 15 15 1 ]
  //: joint g53 (G1) @(362, 175) /w:[ 7 -1 8 14 ]
  and g7 (.I0(Cin), .I1(P0), .I2(G1), .Z(w36));   //: @(536,241) /sn:0 /R:3 /w:[ 11 13 0 1 ]
  and g9 (.I0(Cin), .I1(P0), .Z(w29));   //: @(646,237) /sn:0 /R:3 /w:[ 13 15 0 ]
  //: output g31 (Ps) @(279,366) /sn:0 /R:3 /w:[ 0 ]
  //: input g15 (G0) @(618,98) /sn:0 /R:3 /w:[ 5 ]
  //: input g20 (G3) @(177,92) /sn:0 /R:3 /w:[ 1 ]
  //: joint g39 (P3) @(240, 164) /w:[ 1 -1 2 12 ]
  //: joint g48 (P1) @(402, 180) /w:[ 2 -1 8 1 ]
  //: joint g43 (G1) @(487, 175) /w:[ -1 4 6 3 ]
  //: joint g29 (G0) @(619, 196) /w:[ -1 4 3 6 ]
  //: input g17 (P1) @(505,94) /sn:0 /R:3 /w:[ 5 ]
  //: output g25 (C2) @(380,368) /sn:0 /R:3 /w:[ 0 ]
  //: joint g52 (P1) @(381, 180) /w:[ 9 -1 10 16 ]
  //: joint g42 (G1) @(487, 218) /w:[ 1 2 -1 16 ]
  //: joint g56 (P2) @(245, 187) /w:[ 2 -1 1 18 ]
  and g5 (.I0(G0), .I1(P1), .I2(P2), .Z(w17));   //: @(381,236) /sn:0 /R:3 /w:[ 0 17 11 0 ]
  //: input g14 (P0) @(644,99) /sn:0 /R:3 /w:[ 0 ]
  //: joint g47 (G0) @(510, 196) /w:[ 2 -1 1 8 ]
  //: joint g44 (P2) @(356, 187) /w:[ 6 12 5 14 ]
  //: joint g36 (Cin) @(412, 203) /w:[ 5 -1 6 8 ]
  //: input g21 (P3) @(195,93) /sn:0 /R:3 /w:[ 7 ]
  //: output g24 (C1) @(520,369) /sn:0 /R:3 /w:[ 0 ]
  //: joint g41 (P3) @(215, 164) /w:[ 3 -1 4 10 ]
  //: output g23 (C0) @(621,368) /sn:0 /R:3 /w:[ 0 ]
  //: joint g54 (P2) @(276, 187) /w:[ 4 -1 3 16 ]
  //: joint g40 (P3) @(195, 164) /w:[ 5 6 -1 8 ]
  //: joint g46 (P2) @(376, 187) /w:[ 8 -1 7 10 ]
  //: joint g45 (P1) @(505, 180) /w:[ -1 4 3 6 ]
  //: joint g35 (Gs) @(227, 323) /w:[ -1 2 4 1 ]
  and g0 (.I0(G2), .I1(P3), .Z(w21));   //: @(197,237) /sn:0 /R:3 /w:[ 5 9 1 ]
  //: input g22 (Cin) @(734,203) /sn:0 /R:2 /w:[ 0 ]
  //: output g26 (Gs) @(227,365) /sn:0 /R:3 /w:[ 0 ]
  or g12 (.I0(w36), .I1(w37), .I2(G1), .Z(C1));   //: @(520,292) /sn:0 /R:3 /w:[ 0 0 17 1 ]
  //: input g18 (G2) @(337,92) /sn:0 /R:3 /w:[ 3 ]
  or g33 (.I0(w11), .I1(Gs), .Z(C3));   //: @(84,325) /sn:0 /R:2 /w:[ 1 5 1 ]
  //: joint g30 (P0) @(644, 186) /w:[ -1 1 2 14 ]
  //: joint g49 (P0) @(536, 186) /w:[ 3 -1 4 12 ]

endmodule

module AND(n, p, R, B, A, z);
//: interface  /sz:(40, 40) /bd:[ ]
output p;    //: /sn:0 /dp:1 {0}(652,288)(612,288){1}
output z;    //: /sn:0 /dp:1 {0}(545,331)(548,331)(548,330)(577,330){1}
//: {2}(581,330)(655,330){3}
//: {4}(579,328)(579,290)(591,290){5}
input [15:0] B;    //: /sn:0 {0}(24,426)(63,426){1}
input [15:0] A;    //: /sn:0 {0}(19,245)(65,245){1}
output [15:0] R;    //: /sn:0 /dp:1 {0}(598,197)(358,197)(358,331){1}
//: {2}(360,333)(437,333){3}
//: {4}(356,333)(291,333){5}
output n;    //: /sn:0 /dp:3 {0}(443,258)(514,258){1}
//: {2}(516,256)(516,250)(577,250){3}
//: {4}(581,250)(653,250){5}
//: {6}(579,252)(579,285)(591,285){7}
//: {8}(516,260)(516,294)(524,294){9}
wire w45;    //: /sn:0 {0}(69,391)(149,391){1}
wire w7;    //: /sn:0 {0}(71,220)(148,220){1}
wire w46;    //: /sn:0 {0}(69,381)(149,381){1}
wire w56;    //: /sn:0 {0}(148,300)(71,300){1}
wire w14;    //: /sn:0 {0}(71,270)(148,270){1}
wire w16;    //: /sn:0 {0}(71,250)(148,250){1}
wire w15;    //: /sn:0 {0}(71,260)(148,260){1}
wire w19;    //: /sn:0 {0}(524,359)(508,359)(508,388)(443,388){1}
wire w4;    //: /sn:0 {0}(443,408)(516,408)(516,369)(524,369){1}
wire w38;    //: /sn:0 {0}(69,461)(149,461){1}
wire w3;    //: /sn:0 {0}(71,170)(148,170){1}
wire [15:0] w0;    //: /sn:0 {0}(270,330)(229,330)(229,245)(154,245){1}
wire w37;    //: /sn:0 {0}(69,471)(149,471){1}
wire w34;    //: /sn:0 {0}(71,180)(148,180){1}
wire w43;    //: /sn:0 {0}(69,411)(149,411){1}
wire w21;    //: /sn:0 {0}(443,368)(497,368)(497,349)(524,349){1}
wire [15:0] w58;    //: /sn:0 {0}(155,426)(229,426)(229,335)(270,335){1}
wire w31;    //: /sn:0 {0}(443,268)(513,268)(513,299)(524,299){1}
wire w28;    //: /sn:0 {0}(443,298)(503,298)(503,314)(524,314){1}
wire w36;    //: /sn:0 {0}(69,491)(149,491){1}
wire w41;    //: /sn:0 {0}(69,431)(149,431){1}
wire w20;    //: /sn:0 {0}(443,378)(502,378)(502,354)(524,354){1}
wire w23;    //: /sn:0 {0}(443,348)(489,348)(489,339)(524,339){1}
wire w24;    //: /sn:0 {0}(443,338)(483,338)(483,334)(524,334){1}
wire w1;    //: /sn:0 {0}(71,320)(107,320)(148,320){1}
wire w25;    //: /sn:0 {0}(71,230)(148,230){1}
wire w40;    //: /sn:0 {0}(69,441)(149,441){1}
wire w8;    //: /sn:0 {0}(71,210)(148,210){1}
wire w18;    //: /sn:0 {0}(443,398)(513,398)(513,364)(524,364){1}
wire w30;    //: /sn:0 {0}(443,278)(510,278)(510,304)(524,304){1}
wire w17;    //: /sn:0 {0}(71,240)(148,240){1}
wire w22;    //: /sn:0 {0}(443,358)(493,358)(493,344)(524,344){1}
wire w2;    //: /sn:0 {0}(69,501)(149,501){1}
wire w57;    //: /sn:0 {0}(149,481)(69,481){1}
wire w44;    //: /sn:0 {0}(69,401)(149,401){1}
wire w12;    //: /sn:0 {0}(71,290)(148,290){1}
wire w10;    //: /sn:0 {0}(71,200)(148,200){1}
wire w13;    //: /sn:0 {0}(71,280)(148,280){1}
wire w27;    //: /sn:0 {0}(443,308)(500,308)(500,319)(524,319){1}
wire w48;    //: /sn:0 {0}(69,361)(149,361){1}
wire w5;    //: /sn:0 {0}(71,310)(148,310){1}
wire w33;    //: /sn:0 {0}(71,190)(148,190){1}
wire w47;    //: /sn:0 {0}(69,371)(149,371){1}
wire w29;    //: /sn:0 {0}(443,288)(506,288)(506,309)(524,309){1}
wire w42;    //: /sn:0 {0}(69,421)(149,421){1}
wire w50;    //: /sn:0 {0}(69,351)(149,351){1}
wire w9;    //: /sn:0 {0}(524,329)(483,329)(483,328)(443,328){1}
wire w39;    //: /sn:0 {0}(69,451)(149,451){1}
wire w26;    //: /sn:0 {0}(443,318)(496,318)(496,324)(524,324){1}
//: enddecls

  nor g4 (.I0(n), .I1(z), .Z(p));   //: @(602,288) /sn:0 /w:[ 7 5 1 ]
  //: output g8 (n) @(650,250) /sn:0 /w:[ 5 ]
  //: output g13 (p) @(649,288) /sn:0 /w:[ 0 ]
  //: output g3 (R) @(595,197) /sn:0 /w:[ 0 ]
  and g2 (.I0(w0), .I1(w58), .Z(R));   //: @(281,333) /sn:0 /w:[ 0 1 5 ]
  //: joint g1 (R) @(358, 333) /w:[ 2 1 4 -1 ]
  concat g16 (.I0(w2), .I1(w36), .I2(w57), .I3(w37), .I4(w38), .I5(w39), .I6(w40), .I7(w41), .I8(w42), .I9(w43), .I10(w44), .I11(w45), .I12(w46), .I13(w47), .I14(w48), .I15(w50), .Z(B));   //: @(64,426) /sn:0 /R:2 /w:[ 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:1
  concat g11 (.I0(w4), .I1(w18), .I2(w19), .I3(w20), .I4(w21), .I5(w22), .I6(w23), .I7(w24), .I8(w9), .I9(w26), .I10(w27), .I11(w28), .I12(w29), .I13(w30), .I14(w31), .I15(n), .Z(R));   //: @(438,333) /sn:0 /R:2 /w:[ 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 3 ] /dr:1
  //: joint g6 (n) @(579, 250) /w:[ 4 -1 3 6 ]
  //: joint g9 (z) @(579, 330) /w:[ 2 4 1 -1 ]
  //: input g7 (B) @(22,426) /sn:0 /w:[ 0 ]
  concat g15 (.I0(w1), .I1(w5), .I2(w56), .I3(w12), .I4(w13), .I5(w14), .I6(w15), .I7(w16), .I8(w17), .I9(w25), .I10(w7), .I11(w8), .I12(w10), .I13(w33), .I14(w34), .I15(w3), .Z(A));   //: @(66,245) /sn:0 /R:2 /w:[ 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:1
  concat g17 (.I0(w1), .I1(w5), .I2(w56), .I3(w12), .I4(w13), .I5(w14), .I6(w15), .I7(w16), .I8(w17), .I9(w25), .I10(w7), .I11(w8), .I12(w10), .I13(w33), .I14(w34), .I15(w3), .Z(w0));   //: @(153,245) /sn:0 /w:[ 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 ] /dr:0
  nor g5 (.I0(n), .I1(w31), .I2(w30), .I3(w29), .I4(w28), .I5(w27), .I6(w26), .I7(w9), .I8(w24), .I9(w23), .I10(w22), .I11(w21), .I12(w20), .I13(w19), .I14(w18), .I15(w4), .Z(z));   //: @(535,331) /sn:0 /w:[ 9 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 ]
  //: joint g0 (n) @(516, 258) /w:[ -1 2 1 8 ]
  //: input g22 (A) @(17,245) /sn:0 /w:[ 0 ]
  concat g26 (.I0(w2), .I1(w36), .I2(w57), .I3(w37), .I4(w38), .I5(w39), .I6(w40), .I7(w41), .I8(w42), .I9(w43), .I10(w44), .I11(w45), .I12(w46), .I13(w47), .I14(w48), .I15(w50), .Z(w58));   //: @(154,426) /sn:0 /w:[ 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 ] /dr:0
  //: output g12 (z) @(652,330) /sn:0 /w:[ 3 ]

endmodule
